* NGSPICE file created from test_flat.ext - technology: sky130A

.subckt test_flat clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[0]
+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1]
+ uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
X0 a_25963_4099# a_25759_4581# ua[1].t1 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1 a_24950_4052# bias.Vnbias bias.Vpbias VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.25775 pd=2.41 as=0.145 ps=1.58 w=0.5 l=0.2
X2 a_25963_4672# a_25759_4581# a_25875_4926# VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 VGND.t17 bias.Vnbias a_26985_4099# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=5.08 as=0.6525 ps=5.08 w=2.25 l=0.4
X4 a_25963_4672# a_25759_4581# a_25875_4353# VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X5 VGND.t15 bias.Vnbias a_27540_4099# VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=5.08 as=0.6525 ps=5.08 w=2.25 l=0.4
X6 VGND.t20 a_26430_4353# sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X7 a_25963_4099# a_25759_4581# a_25875_4353# VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X8 VDPWR.t13 bias.Vpbias a_26985_4926# VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
X9 VDPWR.t11 bias.Vpbias a_27540_4926# VDPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
X10 a_24950_4052# a_24690_4014# a_24690_4014# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.17183 pd=1.605 as=0.29 ps=2.58 w=1 l=0.2
X11 ua[1].t0 a_25875_4353# a_25963_4672# VDPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X12 a_26430_4099# a_26430_4353# a_26518_4672# VDPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X13 a_26518_4099# a_25875_4353# a_26430_4099# VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X14 a_25875_4926# a_25875_4353# a_25963_4099# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X15 VGND.t7 a_24690_4014# a_24950_4052# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.17183 ps=1.605 w=1 l=1
X16 bias.Vnbias bias.Vpbias VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.35
X17 a_24690_4014# bias.Vpbias VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
X18 a_26430_4926# a_26430_4353# a_26518_4099# VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X19 a_26518_4672# a_25875_4353# a_26430_4926# VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X20 a_26518_4672# a_25875_4353# a_26430_4353# VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X21 a_26518_4099# a_25875_4353# a_26430_4353# VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X22 a_27073_4099# a_26430_4353# a_26985_4099# VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X23 a_26985_4099# a_25759_4581# a_27073_4672# VDPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X24 a_27540_4099# ua[0].t2 a_27628_4672# VDPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X25 a_27628_4099# a_25759_4581# a_27540_4099# VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X26 VGND.t13 bias.Vnbias bias.Vnbias VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.2
X27 a_26985_4926# a_25759_4581# a_27073_4099# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X28 a_27540_4926# ua[0].t3 a_27628_4099# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.1425 ps=1.285 w=1 l=0.15
X29 VGND.t21 a_25759_4581# sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X30 VGND.t12 bias.Vnbias ua[1].t2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=5.08 as=0.6525 ps=5.08 w=2.25 l=0.4
X31 VGND.t10 bias.Vnbias a_26430_4099# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=5.08 as=0.6525 ps=5.08 w=2.25 l=0.4
X32 a_27073_4672# a_26430_4353# a_26985_4926# VDPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X33 a_27073_4672# a_26430_4353# a_25759_4581# VDPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X34 a_27628_4672# a_25759_4581# a_27540_4926# VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X35 VDPWR.t5 bias.Vpbias a_25875_4926# VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
X36 VDPWR.t3 bias.Vpbias a_26430_4926# VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
X37 a_27628_4672# a_25759_4581# ua[0].t0 VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X38 bias.Vpbias bias.Vpbias VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.35
X39 a_27073_4099# a_26430_4353# a_25759_4581# VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X40 a_27628_4099# a_25759_4581# ua[0].t1 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.1425 pd=1.285 as=0.29 ps=2.58 w=1 l=0.15
X41 VGND.t22 a_25875_4353# sky130_fd_pr__cap_mim_m3_1 l=6 w=3
R0 ua[1].n0 ua[1].t0 449.072
R1 ua[1].n1 ua[1].n0 181.459
R2 ua[1] ua[1].n1 139.065
R3 ua[1].n1 ua[1].t1 132.903
R4 ua[1].n0 ua[1].t2 38.5672
R5 VGND.n20 VGND.n19 18680.8
R6 VGND.n20 VGND.n2 12742.5
R7 VGND.t8 VGND.n20 1969.63
R8 VGND.t5 VGND.n2 604.573
R9 VGND.n12 VGND.n11 590.96
R10 VGND.n19 VGND.n18 590.956
R11 VGND.n16 VGND.n15 590.956
R12 VGND.n14 VGND.n13 590.952
R13 VGND.n22 VGND.n21 394.651
R14 VGND.n1 VGND.t13 230.751
R15 VGND.n15 VGND.t3 215.445
R16 VGND.t18 VGND.n14 215.445
R17 VGND.t1 VGND.n12 215.445
R18 VGND.t0 VGND.t14 213.547
R19 VGND.t16 VGND.t4 213.547
R20 VGND.t9 VGND.t19 213.547
R21 VGND.t11 VGND.t2 213.547
R22 VGND.t6 VGND.t8 170.838
R23 VGND.n21 VGND.t6 120.535
R24 VGND VGND.t7 83.9512
R25 VGND.t3 VGND.t0 82.5717
R26 VGND.t4 VGND.t18 82.5717
R27 VGND.t19 VGND.t1 82.5717
R28 VGND.t2 VGND.t5 82.5717
R29 VGND.n21 VGND.n2 70.2335
R30 VGND.n18 VGND.t15 40.1172
R31 VGND.n11 VGND.t12 40.1172
R32 VGND.n13 VGND.t10 40.1172
R33 VGND.n16 VGND.t17 40.1172
R34 VGND.n6 VGND 18.3754
R35 VGND.n19 VGND.t14 15.186
R36 VGND.n15 VGND.t16 15.186
R37 VGND.n14 VGND.t9 15.186
R38 VGND.n12 VGND.t11 15.186
R39 VGND.n9 VGND.n8 8.22626
R40 VGND.n10 VGND.n9 7.63538
R41 VGND.n18 VGND.n17 6.89244
R42 VGND.n17 VGND.n16 4.54157
R43 VGND.n11 VGND.n10 4.53244
R44 VGND.n13 VGND.n3 4.53244
R45 VGND.n9 VGND.n6 4.12753
R46 VGND.n17 VGND.n3 2.4356
R47 VGND.n10 VGND.n3 2.32017
R48 VGND.n6 VGND.n5 1.8167
R49 VGND.n1 VGND 0.997028
R50 VGND.n4 VGND.t21 0.393176
R51 VGND.n5 VGND.n4 0.327083
R52 VGND VGND.n23 0.269522
R53 VGND.n22 VGND.n1 0.255935
R54 VGND.n23 VGND.n22 0.255935
R55 VGND.n0 VGND 0.236611
R56 VGND.n7 VGND 0.1255
R57 VGND.n23 VGND.n0 0.108139
R58 VGND.n4 VGND.t20 0.0540714
R59 VGND.n5 VGND.t22 0.0540714
R60 VGND.n8 VGND.n0 0.0459545
R61 VGND.n8 VGND.n7 0.0345909
R62 VGND.n7 VGND 0.0175455
R63 VDPWR.n12 VDPWR.t9 651.787
R64 VDPWR.n13 VDPWR.t1 651.431
R65 VDPWR.n2 VDPWR.t10 452.832
R66 VDPWR.n0 VDPWR.t6 434.212
R67 VDPWR.t0 VDPWR.t8 405.264
R68 VDPWR.t10 VDPWR.t19 382.084
R69 VDPWR.t17 VDPWR.t12 382.084
R70 VDPWR.t21 VDPWR.t2 382.084
R71 VDPWR.t4 VDPWR.t15 382.084
R72 VDPWR.n5 VDPWR.n4 379.894
R73 VDPWR.n7 VDPWR.n6 379.892
R74 VDPWR.n9 VDPWR.n8 379.887
R75 VDPWR.n14 VDPWR.n0 379.639
R76 VDPWR.n5 VDPWR.t16 357.771
R77 VDPWR.n7 VDPWR.t20 357.771
R78 VDPWR.n8 VDPWR.t14 357.771
R79 VDPWR.n0 VDPWR.t0 297.368
R80 VDPWR.n4 VDPWR.t13 228.218
R81 VDPWR.n6 VDPWR.t3 228.218
R82 VDPWR.n9 VDPWR.t5 228.218
R83 VDPWR.n2 VDPWR.t11 228.218
R84 VDPWR.n15 VDPWR.t7 228.215
R85 VDPWR.t19 VDPWR.t16 151.097
R86 VDPWR.t20 VDPWR.t17 151.097
R87 VDPWR.t14 VDPWR.t21 151.097
R88 VDPWR.t15 VDPWR.t18 151.097
R89 VDPWR.t12 VDPWR.n5 72.9438
R90 VDPWR.t2 VDPWR.n7 72.9438
R91 VDPWR.n8 VDPWR.t4 72.9438
R92 VDPWR.n11 VDPWR 25.8522
R93 VDPWR.n11 VDPWR.n10 11.3337
R94 VDPWR.n3 VDPWR.n2 6.80678
R95 VDPWR.n12 VDPWR.n11 5.70139
R96 VDPWR.n4 VDPWR.n3 4.5005
R97 VDPWR.n6 VDPWR.n1 4.5005
R98 VDPWR.n10 VDPWR.n9 4.5005
R99 VDPWR.n10 VDPWR.n1 2.36863
R100 VDPWR.n3 VDPWR.n1 2.35524
R101 VDPWR.n15 VDPWR.n14 0.504382
R102 VDPWR.n14 VDPWR.n13 0.371036
R103 VDPWR VDPWR.n15 0.272239
R104 VDPWR.n13 VDPWR.n12 0.13175
R105 ua[0] ua[0].n1 507.483
R106 ua[0].n0 ua[0].t0 278.906
R107 ua[0].n1 ua[0].t2 234.079
R108 ua[0].n1 ua[0].t3 220.484
R109 ua[0].n1 ua[0].n0 202.071
R110 ua[0].n0 ua[0].t1 131.02
C0 a_27628_4099# a_27628_4672# 0.00956f
C1 ua[0] a_25759_4581# 0.409f
C2 a_25875_4926# ua[1] 0.26811f
C3 a_25875_4926# bias.Vnbias 0.0121f
C4 uio_in[1] uio_in[2] 0.03102f
C5 VDPWR a_25759_4581# 0.99799f
C6 uio_out[4] uio_out[3] 0.03102f
C7 a_27540_4926# ua[0] 0.11412f
C8 a_27073_4099# a_25759_4581# 0.2059f
C9 uio_in[1] uio_in[0] 0.03102f
C10 a_26430_4353# a_25759_4581# 1.04813f
C11 a_27540_4926# VDPWR 0.40762f
C12 a_25963_4099# a_25875_4926# 0.16413f
C13 VDPWR a_26430_4099# 0.04811f
C14 uo_out[1] uo_out[2] 0.03102f
C15 ui_in[0] ui_in[1] 0.03102f
C16 a_26430_4353# a_27540_4926# 0.00265f
C17 ui_in[3] ui_in[2] 0.03102f
C18 uio_in[6] uio_in[7] 0.03102f
C19 a_26430_4353# a_26430_4099# 0.18167f
C20 uio_in[4] uio_in[5] 0.03102f
C21 VDPWR ua[0] 0.23806f
C22 ua[1] a_25759_4581# 0.03211f
C23 a_26518_4099# a_26518_4672# 0.00956f
C24 bias.Vnbias a_25759_4581# 0.1344f
C25 uio_oe[0] uio_out[7] 0.03102f
C26 a_24690_4014# a_26518_4099# 0
C27 a_26430_4353# ua[0] 0.00346f
C28 VDPWR a_27073_4099# 0
C29 a_27540_4926# bias.Vnbias 0.00179f
C30 a_26430_4353# VDPWR 0.71702f
C31 a_26430_4099# bias.Vnbias 0.1843f
C32 a_25963_4099# a_25759_4581# 0.02278f
C33 a_26430_4353# a_27073_4099# 0.06693f
C34 a_26430_4926# a_26518_4099# 0.16413f
C35 bias.Vnbias ua[0] 0.01523f
C36 VDPWR ua[1] 0.04849f
C37 uio_out[5] uio_out[6] 0.03102f
C38 VDPWR bias.Vnbias 0.18212f
C39 bias.Vpbias a_27540_4099# 0.00715f
C40 a_27073_4099# bias.Vnbias 0.00138f
C41 a_26430_4353# ua[1] 0.02766f
C42 bias.Vpbias a_26518_4672# 0.03137f
C43 a_26430_4353# bias.Vnbias 0.10982f
C44 a_24690_4014# bias.Vpbias 0.09107f
C45 bias.Vpbias a_26985_4099# 0.00715f
C46 a_25963_4099# VDPWR 0
C47 a_26985_4926# bias.Vpbias 0.11955f
C48 rst_n clk 0.03102f
C49 a_26430_4926# bias.Vpbias 0.12593f
C50 ua[1] bias.Vnbias 0.13708f
C51 a_27628_4672# a_27540_4099# 0.16407f
C52 a_25963_4099# ua[1] 0.26564f
C53 a_25963_4099# bias.Vnbias 0.01485f
C54 a_27073_4672# bias.Vpbias 0.0295f
C55 a_26985_4926# a_27628_4672# 0
C56 a_26518_4672# a_25875_4353# 0.02411f
C57 a_24690_4014# a_25875_4353# 0.01324f
C58 a_26985_4099# a_25875_4353# 0
C59 a_26518_4099# a_25759_4581# 0.01011f
C60 a_26985_4926# a_25875_4353# 0
C61 bias.Vpbias a_25875_4926# 0.16893f
C62 a_26430_4926# a_25875_4353# 0.03876f
C63 a_26518_4099# a_26430_4099# 0.26564f
C64 a_24690_4014# a_24950_4052# 0.01779f
C65 ui_in[2] ui_in[1] 0.03102f
C66 a_26518_4099# VDPWR 0
C67 a_26430_4353# a_26518_4099# 0.21001f
C68 bias.Vpbias a_25759_4581# 0.13408f
C69 a_26430_4926# a_25963_4672# 0.00391f
C70 uio_oe[7] uio_oe[6] 0.03102f
C71 a_27540_4926# bias.Vpbias 0.11844f
C72 uo_out[6] uo_out[5] 0.03102f
C73 bias.Vpbias a_26430_4099# 0.00728f
C74 a_26518_4099# bias.Vnbias 0.00169f
C75 ena clk 0.03102f
C76 a_25875_4926# a_25875_4353# 0.24888f
C77 bias.Vpbias ua[0] 0.01124f
C78 a_27628_4672# a_25759_4581# 0.05368f
C79 a_27628_4099# a_27540_4099# 0.26564f
C80 bias.Vpbias VDPWR 1.24691f
C81 uio_in[4] uio_in[3] 0.03102f
C82 bias.Vpbias a_27073_4099# 0
C83 a_27540_4926# a_27628_4672# 0.28693f
C84 uo_out[7] uio_out[0] 0.03102f
C85 a_26430_4353# bias.Vpbias 0.14459f
C86 a_27628_4672# ua[0] 0.19299f
C87 a_25875_4353# a_25759_4581# 0.55255f
C88 bias.Vpbias ua[1] 0.00786f
C89 a_25875_4926# a_25963_4672# 0.28684f
C90 a_27628_4672# VDPWR 0.06794f
C91 bias.Vpbias bias.Vnbias 0.1915f
C92 a_26430_4099# a_25875_4353# 0.16184f
C93 a_25963_4099# bias.Vpbias 0
C94 uio_out[2] uio_out[1] 0.03102f
C95 a_24950_4052# a_25759_4581# 0
C96 VDPWR a_25875_4353# 0.63859f
C97 a_25963_4672# a_25759_4581# 0.02195f
C98 a_26430_4353# a_25875_4353# 0.63321f
C99 uio_oe[5] uio_oe[4] 0.03102f
C100 uio_in[2] uio_in[3] 0.03102f
C101 uo_out[4] uo_out[5] 0.03102f
C102 ui_in[5] ui_in[6] 0.03102f
C103 a_24950_4052# VDPWR 0.00196f
C104 ua[1] a_25875_4353# 0.23958f
C105 uio_out[0] uio_out[1] 0.03102f
C106 bias.Vnbias a_25875_4353# 0.1626f
C107 VDPWR a_25963_4672# 0.05636f
C108 a_25963_4099# a_25875_4353# 0.23685f
C109 a_27628_4099# a_25759_4581# 0.0712f
C110 a_24950_4052# ua[1] 0
C111 a_24950_4052# bias.Vnbias 0.03669f
C112 a_26985_4926# a_27540_4099# 0
C113 a_27540_4926# a_27628_4099# 0.16413f
C114 a_26985_4926# a_26518_4672# 0.00391f
C115 ua[1] a_25963_4672# 0.16407f
C116 bias.Vnbias a_25963_4672# 0
C117 a_26985_4926# a_26985_4099# 0.26811f
C118 a_26430_4926# a_26518_4672# 0.28684f
C119 ui_in[7] uio_in[0] 0.03102f
C120 a_26430_4926# a_26985_4099# 0
C121 a_27628_4099# ua[0] 0.19568f
C122 a_25963_4099# a_25963_4672# 0.00956f
C123 bias.Vpbias a_26518_4099# 0
C124 uo_out[0] uio_in[7] 0.03102f
C125 a_26985_4926# a_26430_4926# 0.00953f
C126 uio_out[6] uio_out[7] 0.03102f
C127 a_27628_4099# VDPWR 0.0014f
C128 a_27073_4672# a_26985_4099# 0.16407f
C129 a_27073_4672# a_26985_4926# 0.28693f
C130 ui_in[4] ui_in[3] 0.03102f
C131 a_27073_4672# a_26430_4926# 0
C132 a_27628_4099# bias.Vnbias 0.00138f
C133 uio_out[2] uio_out[3] 0.03102f
C134 uio_out[5] uio_out[4] 0.03102f
C135 a_25875_4926# a_26518_4672# 0
C136 a_26518_4099# a_25875_4353# 0.03776f
C137 a_26430_4926# a_25875_4926# 0.00953f
C138 a_27628_4672# bias.Vpbias 0.0295f
C139 uio_oe[4] uio_oe[3] 0.03102f
C140 a_27540_4099# a_25759_4581# 0.26476f
C141 a_26518_4672# a_25759_4581# 0.00929f
C142 a_24690_4014# a_25759_4581# 0
C143 a_26985_4099# a_25759_4581# 0.13245f
C144 a_27540_4926# a_27540_4099# 0.26811f
C145 a_26985_4926# a_25759_4581# 0.17679f
C146 a_26430_4099# a_26518_4672# 0.16407f
C147 ui_in[5] ui_in[4] 0.03102f
C148 a_24690_4014# a_26430_4099# 0
C149 a_26430_4926# a_25759_4581# 0.05777f
C150 bias.Vpbias a_25875_4353# 0.18471f
C151 a_27540_4926# a_26985_4926# 0.00892f
C152 a_27540_4099# ua[0] 0.11412f
C153 uio_oe[1] uio_oe[0] 0.03102f
C154 a_26985_4099# ua[0] 0.02737f
C155 VDPWR a_27540_4099# 0.04951f
C156 a_26430_4926# a_26430_4099# 0.26809f
C157 VDPWR a_26518_4672# 0.06778f
C158 a_26985_4926# ua[0] 0.01388f
C159 a_27073_4672# a_25759_4581# 0.20233f
C160 a_24690_4014# VDPWR 0.14714f
C161 a_26985_4099# VDPWR 0.04814f
C162 uio_oe[5] uio_oe[6] 0.03102f
C163 a_26430_4353# a_27540_4099# 0.00151f
C164 a_26985_4099# a_27073_4099# 0.26564f
C165 a_26430_4353# a_26518_4672# 0.20908f
C166 a_26985_4926# VDPWR 0.40442f
C167 bias.Vpbias a_24950_4052# 0.07529f
C168 uio_oe[3] uio_oe[2] 0.03102f
C169 a_26985_4926# a_27073_4099# 0.16413f
C170 a_26430_4353# a_26985_4099# 0.24146f
C171 a_27073_4672# a_27540_4926# 0.00391f
C172 a_24690_4014# a_26430_4353# 0
C173 a_26430_4926# VDPWR 0.40458f
C174 a_26430_4353# a_26985_4926# 0.12672f
C175 bias.Vpbias a_25963_4672# 0.03951f
C176 ui_in[0] rst_n 0.03102f
C177 a_27540_4099# bias.Vnbias 0.18445f
C178 a_26430_4353# a_26430_4926# 0.20675f
C179 bias.Vnbias a_26518_4672# 0
C180 a_24690_4014# ua[1] 0.00376f
C181 a_24690_4014# bias.Vnbias 0.07372f
C182 a_26985_4099# bias.Vnbias 0.18441f
C183 a_27073_4672# VDPWR 0.06788f
C184 uio_in[6] uio_in[5] 0.03102f
C185 uio_oe[1] uio_oe[2] 0.03102f
C186 a_27073_4672# a_27073_4099# 0.00956f
C187 a_26985_4926# bias.Vnbias 0.00179f
C188 a_25875_4926# a_25759_4581# 0.0623f
C189 a_27073_4672# a_26430_4353# 0.05318f
C190 a_25963_4099# a_24690_4014# 0
C191 a_26430_4926# bias.Vnbias 0.00193f
C192 a_25875_4926# a_26430_4099# 0
C193 uo_out[4] uo_out[3] 0.03102f
C194 uo_out[2] uo_out[3] 0.03102f
C195 uo_out[6] uo_out[7] 0.03102f
C196 ui_in[6] ui_in[7] 0.03102f
C197 a_24950_4052# a_25875_4353# 0.00153f
C198 a_27628_4099# bias.Vpbias 0
C199 uo_out[1] uo_out[0] 0.03102f
C200 a_25875_4926# VDPWR 0.31863f
C201 a_25963_4672# a_25875_4353# 0.23478f
C202 a_26430_4353# a_25875_4926# 0.01422f
C203 a_27540_4926# a_25759_4581# 0.14598f
C204 a_26430_4099# a_25759_4581# 0.04353f
C205 ua[2] VGND 0.14696f
C206 ua[3] VGND 0.14696f
C207 ua[4] VGND 0.14696f
C208 ua[5] VGND 0.14696f
C209 ua[6] VGND 0.14696f
C210 ua[7] VGND 0.14696f
C211 ena VGND 0.07038f
C212 clk VGND 0.04288f
C213 rst_n VGND 0.04288f
C214 ui_in[0] VGND 0.04288f
C215 ui_in[1] VGND 0.04288f
C216 ui_in[2] VGND 0.04288f
C217 ui_in[3] VGND 0.04288f
C218 ui_in[4] VGND 0.04288f
C219 ui_in[5] VGND 0.04288f
C220 ui_in[6] VGND 0.04288f
C221 ui_in[7] VGND 0.04288f
C222 uio_in[0] VGND 0.04288f
C223 uio_in[1] VGND 0.04288f
C224 uio_in[2] VGND 0.04288f
C225 uio_in[3] VGND 0.04288f
C226 uio_in[4] VGND 0.04288f
C227 uio_in[5] VGND 0.04288f
C228 uio_in[6] VGND 0.04288f
C229 uio_in[7] VGND 0.04288f
C230 uo_out[0] VGND 0.04288f
C231 uo_out[1] VGND 0.04288f
C232 uo_out[2] VGND 0.04288f
C233 uo_out[3] VGND 0.04288f
C234 uo_out[4] VGND 0.04288f
C235 uo_out[5] VGND 0.04288f
C236 uo_out[6] VGND 0.04288f
C237 uo_out[7] VGND 0.04288f
C238 uio_out[0] VGND 0.04288f
C239 uio_out[1] VGND 0.04288f
C240 uio_out[2] VGND 0.04288f
C241 uio_out[3] VGND 0.04288f
C242 uio_out[4] VGND 0.04288f
C243 uio_out[5] VGND 0.04288f
C244 uio_out[6] VGND 0.04288f
C245 uio_out[7] VGND 0.04288f
C246 uio_oe[0] VGND 0.04288f
C247 uio_oe[1] VGND 0.04288f
C248 uio_oe[2] VGND 0.04288f
C249 uio_oe[3] VGND 0.04288f
C250 uio_oe[4] VGND 0.04288f
C251 uio_oe[5] VGND 0.04288f
C252 uio_oe[6] VGND 0.04288f
C253 uio_oe[7] VGND 0.07038f
C254 ua[0] VGND 3.86047f
C255 ua[1] VGND 3.09147f
C256 VDPWR VGND 44.2399f
C257 a_27628_4099# VGND 0.08452f
C258 a_27073_4099# VGND 0.08448f
C259 a_26518_4099# VGND 0.09504f
C260 a_25963_4099# VGND 0.08546f
C261 a_24690_4014# VGND 0.8563f
C262 a_24950_4052# VGND 0.07129f
C263 a_27540_4099# VGND 0.56409f
C264 a_27628_4672# VGND 0.02139f
C265 a_26985_4099# VGND 0.52738f
C266 a_27540_4926# VGND 0.18563f
C267 a_27073_4672# VGND 0.01648f
C268 a_26430_4099# VGND 0.54191f
C269 a_26985_4926# VGND 0.15155f
C270 a_26430_4353# VGND 3.5298f
C271 a_26518_4672# VGND 0.02914f
C272 bias.Vnbias VGND 3.07147f
C273 a_26430_4926# VGND 0.16483f
C274 a_25875_4353# VGND 3.86565f
C275 a_25963_4672# VGND 0.01732f
C276 a_25875_4926# VGND 0.19854f
C277 bias.Vpbias VGND 1.80404f
C278 a_25759_4581# VGND 4.47454f
.ends

