magic
tech sky130A
magscale 1 2
timestamp 1738436067
<< checkpaint >>
rect 8 1287 2950 1340
rect 8 1234 3319 1287
rect 8 -2000 3688 1234
rect 377 -2053 3688 -2000
rect 746 -2106 3688 -2053
<< error_s >>
rect 432 987 467 1021
rect 433 968 467 987
rect 241 919 303 925
rect 241 885 253 919
rect 241 879 303 885
rect 241 -409 303 -403
rect 241 -443 253 -409
rect 241 -449 303 -443
rect 452 -545 467 968
rect 486 934 521 968
rect 841 934 876 968
rect 486 -545 520 934
rect 842 915 876 934
rect 650 866 712 872
rect 650 832 662 866
rect 650 826 712 832
rect 650 -462 712 -456
rect 650 -496 662 -462
rect 650 -502 712 -496
rect 486 -579 501 -545
rect 861 -598 876 915
rect 895 881 930 915
rect 895 -598 929 881
rect 1059 813 1121 819
rect 1059 779 1071 813
rect 1059 773 1121 779
rect 1251 80 1285 98
rect 1251 44 1321 80
rect 1268 10 1339 44
rect 1619 10 1654 44
rect 1059 -515 1121 -509
rect 1059 -549 1071 -515
rect 1059 -555 1121 -549
rect 895 -632 910 -598
rect 1268 -651 1338 10
rect 1620 -9 1654 10
rect 1450 -58 1508 -52
rect 1450 -92 1462 -58
rect 1450 -98 1508 -92
rect 1450 -568 1508 -562
rect 1450 -602 1462 -568
rect 1450 -608 1508 -602
rect 1268 -687 1321 -651
rect 1639 -704 1654 -9
rect 1673 -43 1708 -9
rect 1673 -704 1707 -43
rect 1819 -111 1877 -105
rect 1819 -145 1831 -111
rect 1819 -151 1877 -145
rect 1819 -621 1877 -615
rect 1819 -655 1831 -621
rect 1819 -661 1877 -655
rect 1673 -738 1688 -704
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM1
timestamp 1738435636
transform 1 0 1848 0 1 -383
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM2
timestamp 1738435636
transform 1 0 681 0 1 185
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM3
timestamp 1738435636
transform 1 0 2217 0 1 -436
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM4
timestamp 1738435636
transform 1 0 1090 0 1 132
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM6
timestamp 1738435636
transform 1 0 1479 0 1 -330
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM10
timestamp 1738435636
transform 1 0 272 0 1 238
box -231 -819 231 819
<< end >>
