/* Automatically generated from https://wokwi.com/projects/412635532198550529 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_412635532198550529(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = rst_n;
  wire net3 = ui_in[0];
  wire net4 = ui_in[1];
  wire net5 = ui_in[2];
  wire net6 = ui_in[3];
  wire net7 = ui_in[4];
  wire net8 = ui_in[5];
  wire net9 = ui_in[6];
  wire net10 = ui_in[7];
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18;
  wire net19 = uio_in[0];
  wire net20 = 1'b0;
  wire net21 = uio_in[1];
  wire net22 = uio_in[2];
  wire net23 = uio_in[3];
  wire net24 = uio_in[4];
  wire net25 = uio_in[5];
  wire net26;
  wire net27 = 1'b1;
  wire net28;
  wire net29 = 1'b0;
  wire net30 = 1'b1;
  wire net31 = 1'b1;
  wire net32 = 1'b0;
  wire net33 = 1'b1;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103 = 1'b0;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116 = 1'b0;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144 = 1'b1;
  wire net145 = 1'b1;
  wire net146 = 1'b0;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163 = 1'b0;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256 = 1'b0;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265 = 1'b0;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270 = 1'b1;
  wire net271;
  wire net272 = 1'b0;
  wire net273;
  wire net274;
  wire net275;
  wire net276 = 1'b0;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281 = 1'b0;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286 = 1'b0;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291 = 1'b0;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301 = 1'b0;
  wire net302;
  wire net303;
  wire net304 = 1'b0;
  wire net305;
  wire net306;
  wire net307;
  wire net308 = 1'b1;
  wire net309;
  wire net310 = 1'b0;
  wire net311;
  wire net312;
  wire net313;
  wire net314 = 1'b0;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319 = 1'b0;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324 = 1'b0;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329 = 1'b0;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339 = 1'b0;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344 = 1'b0;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349 = 1'b0;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354 = 1'b0;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359 = 1'b0;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369 = 1'b0;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374 = 1'b0;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381 = 1'b0;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386 = 1'b0;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396 = 1'b0;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402 = 1'b0;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428 = 1'b0;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446 = 1'b0;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464 = 1'b0;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;
  wire net474;
  wire net475;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;
  wire net481;
  wire net482 = 1'b0;
  wire net483;
  wire net484;
  wire net485;
  wire net486;
  wire net487;
  wire net488;
  wire net489;
  wire net490;
  wire net491;
  wire net492;
  wire net493;
  wire net494;
  wire net495;
  wire net496;
  wire net497;
  wire net498;
  wire net499;
  wire net500;
  wire net501;
  wire net502;
  wire net503;
  wire net504;
  wire net505;
  wire net506;
  wire net507;
  wire net508;
  wire net509;
  wire net510;
  wire net511;
  wire net512;
  wire net513;
  wire net514;
  wire net515;
  wire net516;
  wire net517;
  wire net518;
  wire net519;
  wire net520;
  wire net521;
  wire net522;
  wire net523;
  wire net524;
  wire net525;
  wire net526;
  wire net527;
  wire net528;
  wire net529;
  wire net530;
  wire net531;
  wire net532;
  wire net533;
  wire net534;
  wire net535;
  wire net536;
  wire net537;
  wire net538;
  wire net539;
  wire net540;
  wire net541;
  wire net542;
  wire net543;
  wire net544;
  wire net545;
  wire net546 = 1'b0;
  wire net547;
  wire net548;
  wire net549;
  wire net550;
  wire net551;
  wire net552;
  wire net553;
  wire net554;
  wire net555;
  wire net556;
  wire net557;
  wire net558;
  wire net559;
  wire net560;
  wire net561;
  wire net562;
  wire net563;
  wire net564;
  wire net565;
  wire net566;
  wire net567;
  wire net568;
  wire net569;
  wire net570 = 1'b1;
  wire net571 = 1'b0;
  wire net572;
  wire net573;
  wire net574;
  wire net575;
  wire net576 = 1'b0;
  wire net577;
  wire net578;
  wire net579;
  wire net580;
  wire net581;
  wire net582;
  wire net583;
  wire net584;
  wire net585;
  wire net586;
  wire net587;
  wire net588;
  wire net589;
  wire net590;
  wire net591;
  wire net592;
  wire net593;
  wire net594;
  wire net595;
  wire net596;
  wire net597;
  wire net598;
  wire net599;
  wire net600;
  wire net601;
  wire net602;
  wire net603;
  wire net604;
  wire net605;
  wire net606;
  wire net607;
  wire net608;
  wire net609;
  wire net610;
  wire net611;
  wire net612;
  wire net613;
  wire net614;
  wire net615;
  wire net616;
  wire net617;
  wire net618;
  wire net619 = 1'b0;
  wire net620;
  wire net621;
  wire net622;
  wire net623;
  wire net624;
  wire net625;
  wire net626;
  wire net627;
  wire net628;
  wire net629;
  wire net630;
  wire net631;
  wire net632;
  wire net633;
  wire net634;
  wire net635;
  wire net636;
  wire net637;
  wire net638;
  wire net639;
  wire net640;
  wire net641;
  wire net642;
  wire net643;
  wire net644;
  wire net645;
  wire net646;
  wire net647;
  wire net648;
  wire net649;
  wire net650;
  wire net651;
  wire net652;
  wire net653;
  wire net654;
  wire net655;
  wire net656;
  wire net657 = 1'b0;
  wire net658 = 1'b0;
  wire net659 = 1'b0;
  wire net660 = 1'b0;
  wire net661;
  wire net662 = 1'b0;
  wire net663;
  wire net664;
  wire net665;
  wire net666 = 1'b0;
  wire net667;
  wire net668;
  wire net669 = 1'b0;
  wire net670;
  wire net671;
  wire net672;
  wire net673;
  wire net674;
  wire net675;
  wire net676;
  wire net677;
  wire net678 = 1'b1;
  wire net679;
  wire net680;
  wire net681;
  wire net682;
  wire net683;
  wire net684;
  wire net685;
  wire net686;
  wire net687;
  wire net688;
  wire net689;
  wire net690;
  wire net691;
  wire net692;
  wire net693;
  wire net694;
  wire net695;
  wire net696;
  wire net697;
  wire net698;
  wire net699;
  wire net700;
  wire net701;
  wire net702;
  wire net703;
  wire net704;
  wire net705 = 1'b0;
  wire net706;
  wire net707;
  wire net708 = 1'b0;
  wire net709 = 1'b0;
  wire net710 = 1'b0;
  wire net711;
  wire net712;
  wire net713;
  wire net714;
  wire net715;
  wire net716;
  wire net717;
  wire net718;

  assign uo_out[0] = net11;
  assign uo_out[1] = net12;
  assign uo_out[2] = net13;
  assign uo_out[3] = net14;
  assign uo_out[4] = net15;
  assign uo_out[5] = net16;
  assign uo_out[6] = net17;
  assign uo_out[7] = net18;
  assign uio_out[0] = net20;
  assign uio_oe[0] = net20;
  assign uio_out[1] = net20;
  assign uio_oe[1] = net20;
  assign uio_out[2] = net20;
  assign uio_oe[2] = net20;
  assign uio_out[3] = net20;
  assign uio_oe[3] = net20;
  assign uio_out[4] = net20;
  assign uio_oe[4] = net20;
  assign uio_out[5] = net20;
  assign uio_oe[5] = net20;
  assign uio_out[6] = net26;
  assign uio_oe[6] = net27;
  assign uio_out[7] = net28;
  assign uio_oe[7] = net27;

  xor_cell xor1 (
    .a (net34),
    .b (net35),
    .out (net36)
  );
  and_cell and1 (
    .a (net37),
    .b (net38),
    .out (net39)
  );
  and_cell and2 (
    .a (net40),
    .b (net37),
    .out (net41)
  );
  and_cell and3 (
    .a (net40),
    .b (net38),
    .out (net42)
  );
  or_cell or3 (
    .a (net39),
    .b (net41),
    .out (net43)
  );
  or_cell or4 (
    .a (net43),
    .b (net42),
    .out (net44)
  );
  and_cell and4 (
    .a (net34),
    .b (net35),
    .out (net45)
  );
  xor_cell xor2 (
    .a (net37),
    .b (net38),
    .out (net46)
  );
  xor_cell xor3 (
    .a (net46),
    .b (net40),
    .out (net47)
  );
  xor_cell xor4 (
    .a (net48),
    .b (net49),
    .out (net50)
  );
  xor_cell xor5 (
    .a (net44),
    .b (net50),
    .out (net51)
  );
  and_cell and5 (
    .a (net48),
    .b (net49),
    .out (net52)
  );
  and_cell and6 (
    .a (net48),
    .b (net44),
    .out (net53)
  );
  and_cell and7 (
    .a (net49),
    .b (net44),
    .out (net54)
  );
  or_cell or1 (
    .a (net52),
    .b (net53),
    .out (net55)
  );
  or_cell or2 (
    .a (net55),
    .b (net54),
    .out (net56)
  );
  xor_cell xor6 (
    .a (net57),
    .b (net58),
    .out (net59)
  );
  xor_cell xor7 (
    .a (net56),
    .b (net59),
    .out (net60)
  );
  and_cell and8 (
    .a (net57),
    .b (net58),
    .out (net61)
  );
  and_cell and9 (
    .a (net57),
    .b (net56),
    .out (net62)
  );
  and_cell and10 (
    .a (net58),
    .b (net56),
    .out (net63)
  );
  or_cell or5 (
    .a (net61),
    .b (net62),
    .out (net64)
  );
  or_cell or6 (
    .a (net64),
    .b (net63),
    .out (net65)
  );
  xor_cell xor8 (
    .a (net66),
    .b (net67),
    .out (net68)
  );
  xor_cell xor9 (
    .a (net65),
    .b (net68),
    .out (net69)
  );
  and_cell and11 (
    .a (net66),
    .b (net67),
    .out (net70)
  );
  and_cell and12 (
    .a (net66),
    .b (net65),
    .out (net71)
  );
  and_cell and13 (
    .a (net67),
    .b (net65),
    .out (net72)
  );
  or_cell or7 (
    .a (net70),
    .b (net71),
    .out (net73)
  );
  or_cell or8 (
    .a (net73),
    .b (net72),
    .out (net74)
  );
  xor_cell xor10 (
    .a (net75),
    .b (net76),
    .out (net77)
  );
  xor_cell xor11 (
    .a (net74),
    .b (net77),
    .out (net78)
  );
  and_cell and14 (
    .a (net75),
    .b (net76),
    .out (net79)
  );
  and_cell and15 (
    .a (net75),
    .b (net74),
    .out (net80)
  );
  and_cell and16 (
    .a (net76),
    .b (net74),
    .out (net81)
  );
  or_cell or9 (
    .a (net79),
    .b (net80),
    .out (net82)
  );
  or_cell or10 (
    .a (net82),
    .b (net81),
    .out (net83)
  );
  xor_cell xor12 (
    .a (net84),
    .b (net85),
    .out (net86)
  );
  xor_cell xor13 (
    .a (net83),
    .b (net86),
    .out (net87)
  );
  and_cell and17 (
    .a (net84),
    .b (net85),
    .out (net88)
  );
  and_cell and18 (
    .a (net84),
    .b (net83),
    .out (net89)
  );
  and_cell and19 (
    .a (net85),
    .b (net83),
    .out (net90)
  );
  or_cell or11 (
    .a (net88),
    .b (net89),
    .out (net91)
  );
  or_cell or12 (
    .a (net91),
    .b (net90),
    .out (net92)
  );
  xor_cell xor14 (
    .a (net93),
    .b (net94),
    .out (net95)
  );
  xor_cell xor15 (
    .a (net92),
    .b (net95),
    .out (net96)
  );
  and_cell and20 (
    .a (net93),
    .b (net94),
    .out (net97)
  );
  and_cell and21 (
    .a (net93),
    .b (net92),
    .out (net98)
  );
  and_cell and22 (
    .a (net94),
    .b (net92),
    .out (net99)
  );
  or_cell or13 (
    .a (net97),
    .b (net98),
    .out (net100)
  );
  or_cell or14 (
    .a (net100),
    .b (net99),
    .out (net101)
  );
  dffsr_cell flop1 (
    .d (net102),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net35),
    .notq ()
  );
  dffsr_cell flop2 (
    .d (net105),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net38),
    .notq ()
  );
  dffsr_cell flop3 (
    .d (net106),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net49),
    .notq ()
  );
  dffsr_cell flop4 (
    .d (net107),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net58),
    .notq ()
  );
  dffsr_cell flop5 (
    .d (net108),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net67),
    .notq ()
  );
  dffsr_cell flop6 (
    .d (net109),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net76),
    .notq ()
  );
  dffsr_cell flop7 (
    .d (net110),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net85),
    .notq ()
  );
  dffsr_cell flop8 (
    .d (net111),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net94),
    .notq ()
  );
  and_cell and24 (
    .a (net112),
    .b (net34),
    .out (net113)
  );
  and_cell and25 (
    .a (net112),
    .b (net35),
    .out (net114)
  );
  or_cell or15 (
    .a (net45),
    .b (net113),
    .out (net115)
  );
  or_cell or16 (
    .a (net115),
    .b (net114),
    .out (net40)
  );
  mux_cell mux1 (
    .a (net116),
    .b (net26),
    .sel (net117),
    .out (net112)
  );
  xor_cell xor16 (
    .a (net36),
    .b (net112),
    .out (net118)
  );
  mux_cell mux2 (
    .a (net119),
    .b (net120),
    .sel (net121),
    .out (net34)
  );
  not_cell not3 (
    .in (net119),
    .out (net122)
  );
  mux_cell mux3 (
    .a (net123),
    .b (net124),
    .sel (net121),
    .out (net37)
  );
  not_cell not4 (
    .in (net123),
    .out (net125)
  );
  mux_cell mux4 (
    .a (net126),
    .b (net127),
    .sel (net121),
    .out (net48)
  );
  not_cell not5 (
    .in (net126),
    .out (net128)
  );
  mux_cell mux5 (
    .a (net129),
    .b (net130),
    .sel (net121),
    .out (net57)
  );
  not_cell not6 (
    .in (net129),
    .out (net131)
  );
  mux_cell mux6 (
    .a (net132),
    .b (net133),
    .sel (net121),
    .out (net66)
  );
  not_cell not7 (
    .in (net132),
    .out (net134)
  );
  mux_cell mux7 (
    .a (net135),
    .b (net136),
    .sel (net121),
    .out (net75)
  );
  not_cell not8 (
    .in (net135),
    .out (net137)
  );
  mux_cell mux8 (
    .a (net138),
    .b (net139),
    .sel (net121),
    .out (net84)
  );
  not_cell not9 (
    .in (net138),
    .out (net140)
  );
  mux_cell mux9 (
    .a (net141),
    .b (net142),
    .sel (net121),
    .out (net93)
  );
  not_cell not10 (
    .in (net141),
    .out (net143)
  );
  dffsr_cell flop9 (
    .d (net21),
    .clk (net1),
    .s (net146),
    .r (net147),
    .q (net148),
    .notq ()
  );
  not_cell not11 (
    .in (net2),
    .out (net147)
  );
  dffsr_cell flop10 (
    .d (net148),
    .clk (net1),
    .s (net146),
    .r (net147),
    .q (net149),
    .notq ()
  );
  dffsr_cell flop11 (
    .d (net149),
    .clk (net1),
    .s (net146),
    .r (net147),
    .q (net150),
    .notq ()
  );
  mux_cell mux10 (
    .a (net151),
    .b (net35),
    .sel (net152),
    .out (net102)
  );
  nand_cell nand1 (
    .a (net153),
    .b (net154),
    .out (net155)
  );
  mux_cell mux11 (
    .a (net156),
    .b (net38),
    .sel (net152),
    .out (net105)
  );
  mux_cell mux12 (
    .a (net157),
    .b (net49),
    .sel (net152),
    .out (net106)
  );
  mux_cell mux13 (
    .a (net158),
    .b (net58),
    .sel (net152),
    .out (net107)
  );
  mux_cell mux14 (
    .a (net159),
    .b (net67),
    .sel (net152),
    .out (net108)
  );
  mux_cell mux15 (
    .a (net160),
    .b (net76),
    .sel (net152),
    .out (net109)
  );
  mux_cell mux16 (
    .a (net161),
    .b (net85),
    .sel (net152),
    .out (net110)
  );
  mux_cell mux17 (
    .a (net162),
    .b (net94),
    .sel (net152),
    .out (net111)
  );
  not_cell not13 (
    .in (net2),
    .out (net104)
  );
  mux_cell mux18 (
    .a (net164),
    .b (net165),
    .sel (net166),
    .out (net167)
  );
  mux_cell mux19 (
    .a (net168),
    .b (net169),
    .sel (net166),
    .out (net170)
  );
  mux_cell mux20 (
    .a (net171),
    .b (net172),
    .sel (net166),
    .out (net173)
  );
  mux_cell mux21 (
    .a (net174),
    .b (net175),
    .sel (net166),
    .out (net176)
  );
  not_cell not14 (
    .in (net167),
    .out (net177)
  );
  not_cell not15 (
    .in (net170),
    .out (net178)
  );
  not_cell not16 (
    .in (net173),
    .out (net179)
  );
  not_cell not17 (
    .in (net176),
    .out (net180)
  );
  and_cell and26 (
    .a (net167),
    .b (net178),
    .out (net181)
  );
  and_cell and27 (
    .a (net181),
    .b (net179),
    .out (net182)
  );
  and_cell and28 (
    .a (net177),
    .b (net170),
    .out (net183)
  );
  and_cell and29 (
    .a (net183),
    .b (net176),
    .out (net184)
  );
  and_cell and30 (
    .a (net178),
    .b (net180),
    .out (net185)
  );
  and_cell and31 (
    .a (net177),
    .b (net173),
    .out (net186)
  );
  and_cell and32 (
    .a (net167),
    .b (net180),
    .out (net187)
  );
  and_cell and33 (
    .a (net170),
    .b (net173),
    .out (net188)
  );
  or_cell or18 (
    .a (net182),
    .b (net184),
    .out (net189)
  );
  or_cell or19 (
    .a (net185),
    .b (net186),
    .out (net190)
  );
  or_cell or20 (
    .a (net187),
    .b (net188),
    .out (net191)
  );
  or_cell or21 (
    .a (net190),
    .b (net191),
    .out (net192)
  );
  or_cell or22 (
    .a (net189),
    .b (net192),
    .out (net193)
  );
  and_cell and34 (
    .a (net177),
    .b (net179),
    .out (net194)
  );
  and_cell and35 (
    .a (net194),
    .b (net180),
    .out (net195)
  );
  and_cell and36 (
    .a (net177),
    .b (net173),
    .out (net196)
  );
  and_cell and37 (
    .a (net196),
    .b (net176),
    .out (net197)
  );
  or_cell or23 (
    .a (net195),
    .b (net197),
    .out (net198)
  );
  and_cell and38 (
    .a (net167),
    .b (net179),
    .out (net199)
  );
  and_cell and39 (
    .a (net199),
    .b (net176),
    .out (net200)
  );
  and_cell and40 (
    .a (net178),
    .b (net179),
    .out (net201)
  );
  and_cell and41 (
    .a (net178),
    .b (net180),
    .out (net202)
  );
  or_cell or24 (
    .a (net201),
    .b (net202),
    .out (net203)
  );
  or_cell or25 (
    .a (net200),
    .b (net203),
    .out (net204)
  );
  or_cell or26 (
    .a (net198),
    .b (net204),
    .out (net205)
  );
  and_cell and42 (
    .a (net177),
    .b (net179),
    .out (net206)
  );
  and_cell and43 (
    .a (net177),
    .b (net176),
    .out (net207)
  );
  and_cell and44 (
    .a (net179),
    .b (net176),
    .out (net208)
  );
  and_cell and45 (
    .a (net177),
    .b (net170),
    .out (net209)
  );
  or_cell or27 (
    .a (net206),
    .b (net207),
    .out (net210)
  );
  or_cell or28 (
    .a (net208),
    .b (net209),
    .out (net211)
  );
  or_cell or29 (
    .a (net210),
    .b (net211),
    .out (net212)
  );
  and_cell and46 (
    .a (net167),
    .b (net178),
    .out (net213)
  );
  or_cell or30 (
    .a (net212),
    .b (net213),
    .out (net214)
  );
  and_cell and47 (
    .a (net177),
    .b (net178),
    .out (net215)
  );
  and_cell and48 (
    .a (net215),
    .b (net180),
    .out (net216)
  );
  and_cell and49 (
    .a (net178),
    .b (net173),
    .out (net217)
  );
  and_cell and50 (
    .a (net217),
    .b (net176),
    .out (net218)
  );
  or_cell or31 (
    .a (net216),
    .b (net218),
    .out (net219)
  );
  and_cell and51 (
    .a (net170),
    .b (net179),
    .out (net220)
  );
  and_cell and52 (
    .a (net220),
    .b (net176),
    .out (net221)
  );
  or_cell or32 (
    .a (net221),
    .b (net222),
    .out (net223)
  );
  or_cell or33 (
    .a (net219),
    .b (net223),
    .out (net224)
  );
  and_cell and53 (
    .a (net170),
    .b (net173),
    .out (net225)
  );
  and_cell and54 (
    .a (net225),
    .b (net180),
    .out (net222)
  );
  and_cell and55 (
    .a (net167),
    .b (net179),
    .out (net226)
  );
  or_cell or34 (
    .a (net224),
    .b (net226),
    .out (net227)
  );
  and_cell and56 (
    .a (net167),
    .b (net173),
    .out (net228)
  );
  and_cell and57 (
    .a (net167),
    .b (net170),
    .out (net229)
  );
  and_cell and58 (
    .a (net173),
    .b (net180),
    .out (net230)
  );
  and_cell and59 (
    .a (net178),
    .b (net180),
    .out (net231)
  );
  or_cell or35 (
    .a (net228),
    .b (net229),
    .out (net232)
  );
  or_cell or36 (
    .a (net230),
    .b (net231),
    .out (net233)
  );
  or_cell or37 (
    .a (net232),
    .b (net233),
    .out (net234)
  );
  and_cell and60 (
    .a (net177),
    .b (net170),
    .out (net235)
  );
  and_cell and61 (
    .a (net235),
    .b (net179),
    .out (net236)
  );
  and_cell and62 (
    .a (net179),
    .b (net180),
    .out (net237)
  );
  and_cell and63 (
    .a (net170),
    .b (net180),
    .out (net238)
  );
  and_cell and64 (
    .a (net167),
    .b (net178),
    .out (net239)
  );
  and_cell and65 (
    .a (net167),
    .b (net173),
    .out (net240)
  );
  or_cell or38 (
    .a (net237),
    .b (net238),
    .out (net241)
  );
  or_cell or39 (
    .a (net239),
    .b (net240),
    .out (net242)
  );
  or_cell or40 (
    .a (net241),
    .b (net242),
    .out (net243)
  );
  or_cell or41 (
    .a (net236),
    .b (net243),
    .out (net244)
  );
  and_cell and66 (
    .a (net177),
    .b (net170),
    .out (net245)
  );
  and_cell and67 (
    .a (net245),
    .b (net179),
    .out (net246)
  );
  and_cell and68 (
    .a (net167),
    .b (net178),
    .out (net247)
  );
  and_cell and69 (
    .a (net167),
    .b (net176),
    .out (net248)
  );
  and_cell and70 (
    .a (net178),
    .b (net173),
    .out (net249)
  );
  and_cell and71 (
    .a (net173),
    .b (net180),
    .out (net250)
  );
  or_cell or42 (
    .a (net247),
    .b (net248),
    .out (net251)
  );
  or_cell or43 (
    .a (net249),
    .b (net250),
    .out (net252)
  );
  or_cell or44 (
    .a (net251),
    .b (net252),
    .out (net253)
  );
  or_cell or45 (
    .a (net246),
    .b (net253),
    .out (net254)
  );
  dffsr_cell flop12 (
    .d (net255),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net11),
    .notq ()
  );
  dffsr_cell flop13 (
    .d (net257),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net12),
    .notq ()
  );
  dffsr_cell flop14 (
    .d (net258),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net13),
    .notq ()
  );
  dffsr_cell flop15 (
    .d (net259),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net14),
    .notq ()
  );
  dffsr_cell flop16 (
    .d (net260),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net15),
    .notq ()
  );
  dffsr_cell flop17 (
    .d (net261),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net16),
    .notq ()
  );
  dffsr_cell flop18 (
    .d (net262),
    .clk (net1),
    .s (net256),
    .r (net104),
    .q (net17),
    .notq ()
  );
  xor_cell xor17 (
    .a (net150),
    .b (net149),
    .out (net263)
  );
  dffsr_cell flop19 (
    .d (net264),
    .clk (net1),
    .s (net265),
    .r (net266),
    .q (net267),
    .notq (net268)
  );
  and_cell and72 (
    .a (net269),
    .b (net147),
    .out (net266)
  );
  not_cell not12 (
    .in (net263),
    .out (net269)
  );
  mux_cell mux22 (
    .a (net267),
    .b (net268),
    .sel (net270),
    .out (net264)
  );
  dffsr_cell flop20 (
    .d (net271),
    .clk (net1),
    .s (net272),
    .r (net266),
    .q (net273),
    .notq (net274)
  );
  mux_cell mux23 (
    .a (net273),
    .b (net274),
    .sel (net267),
    .out (net271)
  );
  dffsr_cell flop21 (
    .d (net275),
    .clk (net1),
    .s (net276),
    .r (net266),
    .q (net277),
    .notq (net278)
  );
  mux_cell mux24 (
    .a (net277),
    .b (net278),
    .sel (net279),
    .out (net275)
  );
  and_cell and74 (
    .a (net273),
    .b (net267),
    .out (net279)
  );
  dffsr_cell flop22 (
    .d (net280),
    .clk (net1),
    .s (net281),
    .r (net266),
    .q (net282),
    .notq (net283)
  );
  mux_cell mux25 (
    .a (net282),
    .b (net283),
    .sel (net284),
    .out (net280)
  );
  and_cell and73 (
    .a (net277),
    .b (net279),
    .out (net284)
  );
  dffsr_cell flop23 (
    .d (net285),
    .clk (net1),
    .s (net286),
    .r (net266),
    .q (net287),
    .notq (net288)
  );
  mux_cell mux26 (
    .a (net287),
    .b (net288),
    .sel (net289),
    .out (net285)
  );
  and_cell and75 (
    .a (net282),
    .b (net284),
    .out (net289)
  );
  dffsr_cell flop24 (
    .d (net290),
    .clk (net1),
    .s (net291),
    .r (net266),
    .q (net292),
    .notq (net293)
  );
  mux_cell mux27 (
    .a (net292),
    .b (net293),
    .sel (net294),
    .out (net290)
  );
  and_cell and76 (
    .a (net287),
    .b (net289),
    .out (net294)
  );
  and_cell and77 (
    .a (net267),
    .b (net273),
    .out (net295)
  );
  and_cell and78 (
    .a (net295),
    .b (net277),
    .out (net296)
  );
  and_cell and79 (
    .a (net296),
    .b (net282),
    .out (net297)
  );
  and_cell and80 (
    .a (net297),
    .b (net287),
    .out (net298)
  );
  and_cell and81 (
    .a (net298),
    .b (net292),
    .out (net299)
  );
  dffsr_cell flop25 (
    .d (net300),
    .clk (net1),
    .s (net301),
    .r (net147),
    .q (net153),
    .notq ()
  );
  mux_cell mux28 (
    .a (net153),
    .b (net149),
    .sel (net299),
    .out (net300)
  );
  dffsr_cell flop26 (
    .d (net153),
    .clk (net1),
    .s (net301),
    .r (net147),
    .q (),
    .notq (net154)
  );
  not_cell not18 (
    .in (net166),
    .out (net302)
  );
  dffsr_cell flop27 (
    .d (net303),
    .clk (net1),
    .s (net304),
    .r (net305),
    .q (net306),
    .notq (net307)
  );
  mux_cell mux29 (
    .a (net306),
    .b (net307),
    .sel (net308),
    .out (net303)
  );
  dffsr_cell flop28 (
    .d (net309),
    .clk (net1),
    .s (net310),
    .r (net305),
    .q (net311),
    .notq (net312)
  );
  mux_cell mux30 (
    .a (net311),
    .b (net312),
    .sel (net306),
    .out (net309)
  );
  dffsr_cell flop29 (
    .d (net313),
    .clk (net1),
    .s (net314),
    .r (net305),
    .q (net315),
    .notq (net316)
  );
  mux_cell mux31 (
    .a (net315),
    .b (net316),
    .sel (net317),
    .out (net313)
  );
  and_cell and83 (
    .a (net311),
    .b (net306),
    .out (net317)
  );
  dffsr_cell flop30 (
    .d (net318),
    .clk (net1),
    .s (net319),
    .r (net305),
    .q (net320),
    .notq (net321)
  );
  mux_cell mux32 (
    .a (net320),
    .b (net321),
    .sel (net322),
    .out (net318)
  );
  and_cell and84 (
    .a (net315),
    .b (net317),
    .out (net322)
  );
  dffsr_cell flop31 (
    .d (net323),
    .clk (net1),
    .s (net324),
    .r (net305),
    .q (net325),
    .notq (net326)
  );
  mux_cell mux33 (
    .a (net325),
    .b (net326),
    .sel (net327),
    .out (net323)
  );
  and_cell and85 (
    .a (net320),
    .b (net322),
    .out (net327)
  );
  dffsr_cell flop32 (
    .d (net328),
    .clk (net1),
    .s (net329),
    .r (net305),
    .q (net330),
    .notq (net331)
  );
  mux_cell mux34 (
    .a (net330),
    .b (net331),
    .sel (net332),
    .out (net328)
  );
  and_cell and86 (
    .a (net325),
    .b (net327),
    .out (net332)
  );
  and_cell and87 (
    .a (net306),
    .b (net311),
    .out (net333)
  );
  and_cell and88 (
    .a (net333),
    .b (net315),
    .out (net334)
  );
  and_cell and89 (
    .a (net334),
    .b (net320),
    .out (net335)
  );
  and_cell and90 (
    .a (net335),
    .b (net325),
    .out (net336)
  );
  and_cell and91 (
    .a (net336),
    .b (net330),
    .out (net337)
  );
  not_cell not19 (
    .in (net2),
    .out (net305)
  );
  dffsr_cell flop33 (
    .d (net338),
    .clk (net1),
    .s (net339),
    .r (net305),
    .q (net340),
    .notq (net341)
  );
  mux_cell mux35 (
    .a (net340),
    .b (net341),
    .sel (net342),
    .out (net338)
  );
  dffsr_cell flop34 (
    .d (net343),
    .clk (net1),
    .s (net344),
    .r (net305),
    .q (net345),
    .notq (net346)
  );
  mux_cell mux36 (
    .a (net345),
    .b (net346),
    .sel (net347),
    .out (net343)
  );
  and_cell and82 (
    .a (net340),
    .b (net342),
    .out (net347)
  );
  dffsr_cell flop35 (
    .d (net348),
    .clk (net1),
    .s (net349),
    .r (net305),
    .q (net350),
    .notq (net351)
  );
  mux_cell mux37 (
    .a (net350),
    .b (net351),
    .sel (net352),
    .out (net348)
  );
  and_cell and92 (
    .a (net345),
    .b (net347),
    .out (net352)
  );
  dffsr_cell flop36 (
    .d (net353),
    .clk (net1),
    .s (net354),
    .r (net305),
    .q (net355),
    .notq (net356)
  );
  mux_cell mux38 (
    .a (net355),
    .b (net356),
    .sel (net357),
    .out (net353)
  );
  and_cell and93 (
    .a (net350),
    .b (net352),
    .out (net357)
  );
  dffsr_cell flop37 (
    .d (net358),
    .clk (net1),
    .s (net359),
    .r (net305),
    .q (net360),
    .notq (net361)
  );
  mux_cell mux39 (
    .a (net360),
    .b (net361),
    .sel (net362),
    .out (net358)
  );
  and_cell and94 (
    .a (net355),
    .b (net357),
    .out (net362)
  );
  and_cell and95 (
    .a (net337),
    .b (net340),
    .out (net363)
  );
  and_cell and96 (
    .a (net363),
    .b (net345),
    .out (net364)
  );
  and_cell and97 (
    .a (net364),
    .b (net350),
    .out (net365)
  );
  and_cell and98 (
    .a (net365),
    .b (net355),
    .out (net366)
  );
  and_cell and99 (
    .a (net366),
    .b (net360),
    .out (net367)
  );
  and_cell and100 (
    .a (net330),
    .b (net332),
    .out (net342)
  );
  dffsr_cell flop38 (
    .d (net368),
    .clk (net1),
    .s (net369),
    .r (net305),
    .q (net370),
    .notq (net371)
  );
  mux_cell mux40 (
    .a (net370),
    .b (net371),
    .sel (net372),
    .out (net368)
  );
  and_cell and101 (
    .a (net360),
    .b (net362),
    .out (net372)
  );
  dffsr_cell flop39 (
    .d (net373),
    .clk (net1),
    .s (net374),
    .r (net305),
    .q (net375),
    .notq (net376)
  );
  mux_cell mux41 (
    .a (net375),
    .b (net376),
    .sel (net377),
    .out (net373)
  );
  and_cell and102 (
    .a (net370),
    .b (net372),
    .out (net377)
  );
  and_cell and103 (
    .a (net367),
    .b (net370),
    .out (net378)
  );
  and_cell and104 (
    .a (net378),
    .b (net375),
    .out (net379)
  );
  dffsr_cell flop40 (
    .d (net380),
    .clk (net1),
    .s (net381),
    .r (net305),
    .q (net382),
    .notq (net383)
  );
  mux_cell mux42 (
    .a (net382),
    .b (net383),
    .sel (net384),
    .out (net380)
  );
  and_cell and105 (
    .a (net375),
    .b (net377),
    .out (net384)
  );
  dffsr_cell flop41 (
    .d (net385),
    .clk (net1),
    .s (net386),
    .r (net305),
    .q (net387),
    .notq (net388)
  );
  mux_cell mux43 (
    .a (net387),
    .b (net388),
    .sel (net389),
    .out (net385)
  );
  and_cell and107 (
    .a (net379),
    .b (net382),
    .out (net390)
  );
  or_cell or46 (
    .a (net391),
    .b (net392),
    .out (net389)
  );
  and_cell and106 (
    .a (net387),
    .b (net393),
    .out (net391)
  );
  and_cell and108 (
    .a (net379),
    .b (net388),
    .out (net392)
  );
  mux_cell mux44 (
    .a (net23),
    .b (net388),
    .sel (net394),
    .out (net166)
  );
  dffsr_cell flop42 (
    .d (net395),
    .clk (net1),
    .s (net396),
    .r (net305),
    .q (net397),
    .notq (net398)
  );
  mux_cell mux45 (
    .a (net397),
    .b (net398),
    .sel (net399),
    .out (net395)
  );
  and_cell and109 (
    .a (net382),
    .b (net384),
    .out (net399)
  );
  and_cell and110 (
    .a (net390),
    .b (net397),
    .out (net393)
  );
  mux_cell mux46 (
    .a (net118),
    .b (net34),
    .sel (net400),
    .out (net151)
  );
  mux_cell mux47 (
    .a (net47),
    .b (net37),
    .sel (net400),
    .out (net156)
  );
  mux_cell mux48 (
    .a (net51),
    .b (net48),
    .sel (net400),
    .out (net157)
  );
  mux_cell mux49 (
    .a (net60),
    .b (net57),
    .sel (net400),
    .out (net158)
  );
  mux_cell mux50 (
    .a (net69),
    .b (net66),
    .sel (net400),
    .out (net159)
  );
  mux_cell mux51 (
    .a (net78),
    .b (net75),
    .sel (net400),
    .out (net160)
  );
  mux_cell mux52 (
    .a (net87),
    .b (net84),
    .sel (net400),
    .out (net161)
  );
  mux_cell mux53 (
    .a (net96),
    .b (net93),
    .sel (net400),
    .out (net162)
  );
  dffsr_cell flop43 (
    .d (net401),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net403),
    .notq ()
  );
  dffsr_cell flop44 (
    .d (net404),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net405),
    .notq ()
  );
  dffsr_cell flop45 (
    .d (net406),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net407),
    .notq ()
  );
  dffsr_cell flop46 (
    .d (net408),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net409),
    .notq ()
  );
  dffsr_cell flop47 (
    .d (net410),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net411),
    .notq ()
  );
  dffsr_cell flop48 (
    .d (net412),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net413),
    .notq ()
  );
  dffsr_cell flop49 (
    .d (net414),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net415),
    .notq ()
  );
  dffsr_cell flop50 (
    .d (net416),
    .clk (net1),
    .s (net402),
    .r (net305),
    .q (net417),
    .notq ()
  );
  mux_cell mux54 (
    .a (net418),
    .b (net403),
    .sel (net419),
    .out (net401)
  );
  mux_cell mux55 (
    .a (net420),
    .b (net405),
    .sel (net419),
    .out (net404)
  );
  mux_cell mux56 (
    .a (net421),
    .b (net407),
    .sel (net419),
    .out (net406)
  );
  mux_cell mux57 (
    .a (net422),
    .b (net409),
    .sel (net419),
    .out (net408)
  );
  mux_cell mux58 (
    .a (net423),
    .b (net411),
    .sel (net419),
    .out (net410)
  );
  mux_cell mux59 (
    .a (net424),
    .b (net413),
    .sel (net419),
    .out (net412)
  );
  mux_cell mux60 (
    .a (net425),
    .b (net415),
    .sel (net419),
    .out (net414)
  );
  mux_cell mux61 (
    .a (net426),
    .b (net417),
    .sel (net419),
    .out (net416)
  );
  dffsr_cell flop51 (
    .d (net427),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net429),
    .notq ()
  );
  dffsr_cell flop52 (
    .d (net430),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net431),
    .notq ()
  );
  dffsr_cell flop53 (
    .d (net432),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net433),
    .notq ()
  );
  dffsr_cell flop54 (
    .d (net434),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net435),
    .notq ()
  );
  dffsr_cell flop55 (
    .d (net436),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net437),
    .notq ()
  );
  dffsr_cell flop56 (
    .d (net438),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net439),
    .notq ()
  );
  dffsr_cell flop57 (
    .d (net440),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net441),
    .notq ()
  );
  dffsr_cell flop58 (
    .d (net442),
    .clk (net1),
    .s (net428),
    .r (net305),
    .q (net443),
    .notq ()
  );
  mux_cell mux62 (
    .a (net418),
    .b (net429),
    .sel (net444),
    .out (net427)
  );
  mux_cell mux63 (
    .a (net420),
    .b (net431),
    .sel (net444),
    .out (net430)
  );
  mux_cell mux64 (
    .a (net421),
    .b (net433),
    .sel (net444),
    .out (net432)
  );
  mux_cell mux65 (
    .a (net422),
    .b (net435),
    .sel (net444),
    .out (net434)
  );
  mux_cell mux66 (
    .a (net423),
    .b (net437),
    .sel (net444),
    .out (net436)
  );
  mux_cell mux67 (
    .a (net424),
    .b (net439),
    .sel (net444),
    .out (net438)
  );
  mux_cell mux68 (
    .a (net425),
    .b (net441),
    .sel (net444),
    .out (net440)
  );
  mux_cell mux69 (
    .a (net426),
    .b (net443),
    .sel (net444),
    .out (net442)
  );
  dffsr_cell flop59 (
    .d (net445),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net447),
    .notq ()
  );
  dffsr_cell flop60 (
    .d (net448),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net449),
    .notq ()
  );
  dffsr_cell flop61 (
    .d (net450),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net451),
    .notq ()
  );
  dffsr_cell flop62 (
    .d (net452),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net453),
    .notq ()
  );
  dffsr_cell flop63 (
    .d (net454),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net455),
    .notq ()
  );
  dffsr_cell flop64 (
    .d (net456),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net457),
    .notq ()
  );
  dffsr_cell flop65 (
    .d (net458),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net459),
    .notq ()
  );
  dffsr_cell flop66 (
    .d (net460),
    .clk (net1),
    .s (net446),
    .r (net305),
    .q (net461),
    .notq ()
  );
  mux_cell mux70 (
    .a (net418),
    .b (net447),
    .sel (net462),
    .out (net445)
  );
  mux_cell mux71 (
    .a (net420),
    .b (net449),
    .sel (net462),
    .out (net448)
  );
  mux_cell mux72 (
    .a (net421),
    .b (net451),
    .sel (net462),
    .out (net450)
  );
  mux_cell mux73 (
    .a (net422),
    .b (net453),
    .sel (net462),
    .out (net452)
  );
  mux_cell mux74 (
    .a (net423),
    .b (net455),
    .sel (net462),
    .out (net454)
  );
  mux_cell mux75 (
    .a (net424),
    .b (net457),
    .sel (net462),
    .out (net456)
  );
  mux_cell mux76 (
    .a (net425),
    .b (net459),
    .sel (net462),
    .out (net458)
  );
  mux_cell mux77 (
    .a (net426),
    .b (net461),
    .sel (net462),
    .out (net460)
  );
  dffsr_cell flop67 (
    .d (net463),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net465),
    .notq ()
  );
  dffsr_cell flop68 (
    .d (net466),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net467),
    .notq ()
  );
  dffsr_cell flop69 (
    .d (net468),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net469),
    .notq ()
  );
  dffsr_cell flop70 (
    .d (net470),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net471),
    .notq ()
  );
  dffsr_cell flop71 (
    .d (net472),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net473),
    .notq ()
  );
  dffsr_cell flop72 (
    .d (net474),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net475),
    .notq ()
  );
  dffsr_cell flop73 (
    .d (net476),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net477),
    .notq ()
  );
  dffsr_cell flop74 (
    .d (net478),
    .clk (net1),
    .s (net464),
    .r (net305),
    .q (net479),
    .notq ()
  );
  mux_cell mux78 (
    .a (net418),
    .b (net465),
    .sel (net480),
    .out (net463)
  );
  mux_cell mux79 (
    .a (net420),
    .b (net467),
    .sel (net480),
    .out (net466)
  );
  mux_cell mux80 (
    .a (net421),
    .b (net469),
    .sel (net480),
    .out (net468)
  );
  mux_cell mux81 (
    .a (net422),
    .b (net471),
    .sel (net480),
    .out (net470)
  );
  mux_cell mux82 (
    .a (net423),
    .b (net473),
    .sel (net480),
    .out (net472)
  );
  mux_cell mux83 (
    .a (net424),
    .b (net475),
    .sel (net480),
    .out (net474)
  );
  mux_cell mux84 (
    .a (net425),
    .b (net477),
    .sel (net480),
    .out (net476)
  );
  mux_cell mux85 (
    .a (net426),
    .b (net479),
    .sel (net480),
    .out (net478)
  );
  mux_cell mux86 (
    .a (net481),
    .b (net481),
    .sel (net482),
    .out (net483)
  );
  mux_cell mux87 (
    .a (net484),
    .b (net484),
    .sel (net482),
    .out (net485)
  );
  not_cell not1 (
    .in (net485),
    .out (net486)
  );
  not_cell not2 (
    .in (net483),
    .out (net487)
  );
  and_cell and111 (
    .a (net487),
    .b (net486),
    .out (net488)
  );
  and_cell and113 (
    .a (net483),
    .b (net486),
    .out (net489)
  );
  and_cell and115 (
    .a (net487),
    .b (net485),
    .out (net490)
  );
  and_cell and117 (
    .a (net483),
    .b (net485),
    .out (net491)
  );
  mux_cell mux88 (
    .a (net151),
    .b (net35),
    .sel (net492),
    .out (net418)
  );
  mux_cell mux89 (
    .a (net156),
    .b (net38),
    .sel (net492),
    .out (net420)
  );
  mux_cell mux90 (
    .a (net157),
    .b (net49),
    .sel (net492),
    .out (net421)
  );
  mux_cell mux91 (
    .a (net158),
    .b (net58),
    .sel (net492),
    .out (net422)
  );
  mux_cell mux92 (
    .a (net159),
    .b (net67),
    .sel (net492),
    .out (net423)
  );
  mux_cell mux93 (
    .a (net160),
    .b (net76),
    .sel (net492),
    .out (net424)
  );
  mux_cell mux94 (
    .a (net161),
    .b (net85),
    .sel (net492),
    .out (net425)
  );
  mux_cell mux95 (
    .a (net162),
    .b (net94),
    .sel (net492),
    .out (net426)
  );
  mux_cell mux96 (
    .a (net429),
    .b (net403),
    .sel (net493),
    .out (net494)
  );
  mux_cell mux97 (
    .a (net431),
    .b (net405),
    .sel (net493),
    .out (net495)
  );
  mux_cell mux98 (
    .a (net433),
    .b (net407),
    .sel (net493),
    .out (net496)
  );
  mux_cell mux99 (
    .a (net435),
    .b (net409),
    .sel (net493),
    .out (net497)
  );
  mux_cell mux100 (
    .a (net437),
    .b (net411),
    .sel (net493),
    .out (net498)
  );
  mux_cell mux101 (
    .a (net439),
    .b (net413),
    .sel (net493),
    .out (net499)
  );
  mux_cell mux102 (
    .a (net441),
    .b (net415),
    .sel (net493),
    .out (net500)
  );
  mux_cell mux103 (
    .a (net443),
    .b (net417),
    .sel (net493),
    .out (net501)
  );
  mux_cell mux104 (
    .a (net465),
    .b (net447),
    .sel (net493),
    .out (net502)
  );
  mux_cell mux105 (
    .a (net467),
    .b (net449),
    .sel (net493),
    .out (net503)
  );
  mux_cell mux106 (
    .a (net469),
    .b (net451),
    .sel (net493),
    .out (net504)
  );
  mux_cell mux107 (
    .a (net471),
    .b (net453),
    .sel (net493),
    .out (net505)
  );
  mux_cell mux108 (
    .a (net473),
    .b (net455),
    .sel (net493),
    .out (net506)
  );
  mux_cell mux109 (
    .a (net475),
    .b (net457),
    .sel (net493),
    .out (net507)
  );
  mux_cell mux110 (
    .a (net477),
    .b (net459),
    .sel (net493),
    .out (net508)
  );
  mux_cell mux111 (
    .a (net479),
    .b (net461),
    .sel (net493),
    .out (net509)
  );
  mux_cell mux112 (
    .a (net502),
    .b (net494),
    .sel (net510),
    .out (net511)
  );
  mux_cell mux113 (
    .a (net503),
    .b (net495),
    .sel (net510),
    .out (net512)
  );
  mux_cell mux114 (
    .a (net504),
    .b (net496),
    .sel (net510),
    .out (net513)
  );
  mux_cell mux115 (
    .a (net505),
    .b (net497),
    .sel (net510),
    .out (net514)
  );
  mux_cell mux116 (
    .a (net506),
    .b (net498),
    .sel (net510),
    .out (net515)
  );
  mux_cell mux117 (
    .a (net507),
    .b (net499),
    .sel (net510),
    .out (net516)
  );
  mux_cell mux118 (
    .a (net508),
    .b (net500),
    .sel (net510),
    .out (net517)
  );
  mux_cell mux119 (
    .a (net509),
    .b (net501),
    .sel (net510),
    .out (net518)
  );
  mux_cell mux120 (
    .a (net519),
    .b (net3),
    .sel (net520),
    .out (net119)
  );
  mux_cell mux121 (
    .a (net521),
    .b (net4),
    .sel (net520),
    .out (net123)
  );
  mux_cell mux122 (
    .a (net522),
    .b (net5),
    .sel (net520),
    .out (net126)
  );
  mux_cell mux123 (
    .a (net523),
    .b (net6),
    .sel (net520),
    .out (net129)
  );
  mux_cell mux124 (
    .a (net524),
    .b (net8),
    .sel (net520),
    .out (net135)
  );
  mux_cell mux125 (
    .a (net525),
    .b (net7),
    .sel (net520),
    .out (net132)
  );
  mux_cell mux126 (
    .a (net526),
    .b (net9),
    .sel (net520),
    .out (net138)
  );
  mux_cell mux127 (
    .a (net527),
    .b (net10),
    .sel (net520),
    .out (net141)
  );
  mux_cell mux128 (
    .a (net528),
    .b (net529),
    .sel (net530),
    .out (net519)
  );
  mux_cell mux129 (
    .a (net531),
    .b (net532),
    .sel (net530),
    .out (net521)
  );
  mux_cell mux130 (
    .a (net533),
    .b (net534),
    .sel (net530),
    .out (net522)
  );
  mux_cell mux131 (
    .a (net535),
    .b (net536),
    .sel (net530),
    .out (net523)
  );
  mux_cell mux132 (
    .a (net537),
    .b (net538),
    .sel (net530),
    .out (net525)
  );
  mux_cell mux133 (
    .a (net539),
    .b (net540),
    .sel (net530),
    .out (net524)
  );
  mux_cell mux134 (
    .a (net541),
    .b (net542),
    .sel (net530),
    .out (net526)
  );
  mux_cell mux135 (
    .a (net543),
    .b (net544),
    .sel (net530),
    .out (net527)
  );
  dffsr_cell flop75 (
    .d (net545),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net481),
    .notq (net548)
  );
  dffsr_cell flop76 (
    .d (net549),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net484),
    .notq (net550)
  );
  dffsr_cell flop77 (
    .d (net551),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net552),
    .notq (net553)
  );
  dffsr_cell flop78 (
    .d (net554),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net555),
    .notq (net556)
  );
  dffsr_cell flop79 (
    .d (net557),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net558),
    .notq (net559)
  );
  dffsr_cell flop80 (
    .d (net560),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net561),
    .notq (net520)
  );
  dffsr_cell flop81 (
    .d (net562),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net400),
    .notq (net563)
  );
  dffsr_cell flop82 (
    .d (net564),
    .clk (net1),
    .s (net546),
    .r (net547),
    .q (net565),
    .notq (net566)
  );
  mux_cell mux136 (
    .a (net3),
    .b (net481),
    .sel (net567),
    .out (net545)
  );
  mux_cell mux137 (
    .a (net4),
    .b (net484),
    .sel (net567),
    .out (net549)
  );
  mux_cell mux138 (
    .a (net5),
    .b (net552),
    .sel (net567),
    .out (net551)
  );
  mux_cell mux139 (
    .a (net6),
    .b (net555),
    .sel (net567),
    .out (net554)
  );
  mux_cell mux140 (
    .a (net7),
    .b (net558),
    .sel (net567),
    .out (net557)
  );
  mux_cell mux141 (
    .a (net8),
    .b (net561),
    .sel (net567),
    .out (net560)
  );
  mux_cell mux142 (
    .a (net9),
    .b (net400),
    .sel (net567),
    .out (net562)
  );
  mux_cell mux143 (
    .a (net10),
    .b (net565),
    .sel (net567),
    .out (net564)
  );
  not_cell not20 (
    .in (net2),
    .out (net547)
  );
  and_cell and118 (
    .a (net565),
    .b (net568),
    .out (net569)
  );
  and_cell and120 (
    .a (net558),
    .b (net563),
    .out (net121)
  );
  not_cell not22 (
    .in (net19),
    .out (net567)
  );
  or_cell or17 (
    .a (net572),
    .b (net155),
    .out (net152)
  );
  nand_cell nand2 (
    .a (net488),
    .b (net569),
    .out (net419)
  );
  not_cell not21 (
    .in (net155),
    .out (net568)
  );
  nand_cell nand3 (
    .a (net489),
    .b (net569),
    .out (net444)
  );
  nand_cell nand4 (
    .a (net490),
    .b (net569),
    .out (net462)
  );
  nand_cell nand5 (
    .a (net491),
    .b (net569),
    .out (net480)
  );
  and_cell and23 (
    .a (net400),
    .b (net565),
    .out (net573)
  );
  and_cell and112 (
    .a (net558),
    .b (net520),
    .out (net574)
  );
  and_cell and114 (
    .a (net574),
    .b (net573),
    .out (net492)
  );
  mux_cell mux144 (
    .a (net193),
    .b (net174),
    .sel (net22),
    .out (net255)
  );
  mux_cell mux145 (
    .a (net205),
    .b (net171),
    .sel (net22),
    .out (net257)
  );
  mux_cell mux146 (
    .a (net214),
    .b (net168),
    .sel (net22),
    .out (net258)
  );
  mux_cell mux147 (
    .a (net227),
    .b (net164),
    .sel (net22),
    .out (net259)
  );
  mux_cell mux148 (
    .a (net234),
    .b (net175),
    .sel (net22),
    .out (net260)
  );
  mux_cell mux149 (
    .a (net244),
    .b (net172),
    .sel (net22),
    .out (net261)
  );
  mux_cell mux150 (
    .a (net254),
    .b (net169),
    .sel (net22),
    .out (net262)
  );
  not_cell not23 (
    .in (net24),
    .out (net394)
  );
  dffsr_cell flop83 (
    .d (net575),
    .clk (net1),
    .s (net576),
    .r (net104),
    .q (net18),
    .notq ()
  );
  mux_cell mux151 (
    .a (net302),
    .b (net165),
    .sel (net22),
    .out (net575)
  );
  mux_cell mux152 (
    .a (net49),
    .b (net157),
    .sel (net25),
    .out (net168)
  );
  mux_cell mux153 (
    .a (net58),
    .b (net158),
    .sel (net25),
    .out (net164)
  );
  mux_cell mux154 (
    .a (net67),
    .b (net159),
    .sel (net25),
    .out (net175)
  );
  mux_cell mux155 (
    .a (net76),
    .b (net160),
    .sel (net25),
    .out (net172)
  );
  mux_cell mux156 (
    .a (net85),
    .b (net161),
    .sel (net25),
    .out (net169)
  );
  mux_cell mux157 (
    .a (net38),
    .b (net156),
    .sel (net25),
    .out (net171)
  );
  mux_cell mux158 (
    .a (net35),
    .b (net151),
    .sel (net25),
    .out (net174)
  );
  mux_cell mux159 (
    .a (net94),
    .b (net162),
    .sel (net25),
    .out (net165)
  );
  and_cell and119 (
    .a (net561),
    .b (net565),
    .out (net577)
  );
  mux_cell mux160 (
    .a (net550),
    .b (net556),
    .sel (net577),
    .out (net510)
  );
  mux_cell mux161 (
    .a (net548),
    .b (net553),
    .sel (net577),
    .out (net493)
  );
  and_cell and116 (
    .a (net35),
    .b (net511),
    .out (net578)
  );
  and_cell and121 (
    .a (net38),
    .b (net512),
    .out (net579)
  );
  and_cell and122 (
    .a (net49),
    .b (net513),
    .out (net580)
  );
  and_cell and123 (
    .a (net58),
    .b (net514),
    .out (net581)
  );
  and_cell and124 (
    .a (net67),
    .b (net515),
    .out (net582)
  );
  and_cell and125 (
    .a (net76),
    .b (net516),
    .out (net583)
  );
  and_cell and126 (
    .a (net85),
    .b (net517),
    .out (net584)
  );
  and_cell and127 (
    .a (net94),
    .b (net518),
    .out (net585)
  );
  or_cell or47 (
    .a (net35),
    .b (net511),
    .out (net586)
  );
  or_cell or48 (
    .a (net38),
    .b (net512),
    .out (net587)
  );
  or_cell or49 (
    .a (net49),
    .b (net513),
    .out (net588)
  );
  or_cell or50 (
    .a (net58),
    .b (net514),
    .out (net589)
  );
  or_cell or51 (
    .a (net67),
    .b (net515),
    .out (net590)
  );
  or_cell or52 (
    .a (net76),
    .b (net516),
    .out (net591)
  );
  or_cell or53 (
    .a (net85),
    .b (net517),
    .out (net592)
  );
  or_cell or54 (
    .a (net94),
    .b (net518),
    .out (net593)
  );
  xor_cell xor18 (
    .a (net35),
    .b (net511),
    .out (net594)
  );
  xor_cell xor19 (
    .a (net38),
    .b (net512),
    .out (net595)
  );
  xor_cell xor20 (
    .a (net49),
    .b (net513),
    .out (net596)
  );
  xor_cell xor21 (
    .a (net58),
    .b (net514),
    .out (net597)
  );
  xor_cell xor22 (
    .a (net67),
    .b (net515),
    .out (net598)
  );
  xor_cell xor23 (
    .a (net76),
    .b (net516),
    .out (net599)
  );
  xor_cell xor24 (
    .a (net85),
    .b (net517),
    .out (net600)
  );
  xor_cell xor25 (
    .a (net94),
    .b (net518),
    .out (net601)
  );
  mux_cell mux162 (
    .a (net586),
    .b (net578),
    .sel (net602),
    .out (net603)
  );
  mux_cell mux163 (
    .a (net587),
    .b (net579),
    .sel (net602),
    .out (net604)
  );
  mux_cell mux164 (
    .a (net588),
    .b (net580),
    .sel (net602),
    .out (net605)
  );
  mux_cell mux165 (
    .a (net589),
    .b (net581),
    .sel (net602),
    .out (net606)
  );
  mux_cell mux166 (
    .a (net590),
    .b (net582),
    .sel (net602),
    .out (net607)
  );
  mux_cell mux167 (
    .a (net591),
    .b (net583),
    .sel (net602),
    .out (net608)
  );
  mux_cell mux168 (
    .a (net592),
    .b (net584),
    .sel (net602),
    .out (net609)
  );
  mux_cell mux169 (
    .a (net593),
    .b (net585),
    .sel (net602),
    .out (net610)
  );
  mux_cell mux170 (
    .a (net511),
    .b (net594),
    .sel (net602),
    .out (net611)
  );
  mux_cell mux171 (
    .a (net512),
    .b (net595),
    .sel (net602),
    .out (net612)
  );
  mux_cell mux172 (
    .a (net513),
    .b (net596),
    .sel (net602),
    .out (net613)
  );
  mux_cell mux173 (
    .a (net514),
    .b (net597),
    .sel (net602),
    .out (net614)
  );
  mux_cell mux174 (
    .a (net515),
    .b (net598),
    .sel (net602),
    .out (net615)
  );
  mux_cell mux175 (
    .a (net516),
    .b (net599),
    .sel (net602),
    .out (net616)
  );
  mux_cell mux176 (
    .a (net517),
    .b (net600),
    .sel (net602),
    .out (net617)
  );
  mux_cell mux177 (
    .a (net518),
    .b (net601),
    .sel (net602),
    .out (net618)
  );
  not_cell not24 (
    .in (net35),
    .out (net620)
  );
  not_cell not25 (
    .in (net38),
    .out (net621)
  );
  not_cell not26 (
    .in (net49),
    .out (net622)
  );
  not_cell not27 (
    .in (net58),
    .out (net623)
  );
  not_cell not28 (
    .in (net67),
    .out (net624)
  );
  not_cell not29 (
    .in (net76),
    .out (net625)
  );
  not_cell not30 (
    .in (net85),
    .out (net626)
  );
  not_cell not31 (
    .in (net94),
    .out (net627)
  );
  not_cell not32 (
    .in (net511),
    .out (net628)
  );
  not_cell not33 (
    .in (net512),
    .out (net629)
  );
  not_cell not34 (
    .in (net513),
    .out (net630)
  );
  not_cell not35 (
    .in (net514),
    .out (net631)
  );
  not_cell not36 (
    .in (net515),
    .out (net632)
  );
  not_cell not37 (
    .in (net516),
    .out (net633)
  );
  not_cell not38 (
    .in (net517),
    .out (net634)
  );
  not_cell not39 (
    .in (net518),
    .out (net635)
  );
  and_cell and128 (
    .a (net636),
    .b (net552),
    .out (net602)
  );
  mux_cell mux178 (
    .a (net628),
    .b (net637),
    .sel (net553),
    .out (net638)
  );
  mux_cell mux179 (
    .a (net629),
    .b (net639),
    .sel (net553),
    .out (net640)
  );
  mux_cell mux180 (
    .a (net630),
    .b (net641),
    .sel (net553),
    .out (net642)
  );
  mux_cell mux181 (
    .a (net631),
    .b (net643),
    .sel (net553),
    .out (net644)
  );
  mux_cell mux182 (
    .a (net632),
    .b (net645),
    .sel (net553),
    .out (net646)
  );
  mux_cell mux183 (
    .a (net633),
    .b (net647),
    .sel (net553),
    .out (net648)
  );
  mux_cell mux184 (
    .a (net634),
    .b (net649),
    .sel (net553),
    .out (net650)
  );
  mux_cell mux185 (
    .a (net635),
    .b (net651),
    .sel (net553),
    .out (net652)
  );
  mux_cell mux186 (
    .a (net611),
    .b (net603),
    .sel (net653),
    .out (net528)
  );
  mux_cell mux187 (
    .a (net612),
    .b (net604),
    .sel (net653),
    .out (net531)
  );
  mux_cell mux188 (
    .a (net613),
    .b (net605),
    .sel (net653),
    .out (net533)
  );
  mux_cell mux189 (
    .a (net614),
    .b (net606),
    .sel (net653),
    .out (net535)
  );
  mux_cell mux190 (
    .a (net615),
    .b (net607),
    .sel (net653),
    .out (net537)
  );
  mux_cell mux191 (
    .a (net616),
    .b (net608),
    .sel (net653),
    .out (net539)
  );
  mux_cell mux192 (
    .a (net617),
    .b (net609),
    .sel (net653),
    .out (net541)
  );
  mux_cell mux193 (
    .a (net618),
    .b (net610),
    .sel (net653),
    .out (net543)
  );
  and_cell and129 (
    .a (net400),
    .b (net566),
    .out (net654)
  );
  and_cell and130 (
    .a (net559),
    .b (net561),
    .out (net655)
  );
  and_cell and131 (
    .a (net636),
    .b (net555),
    .out (net653)
  );
  and_cell and132 (
    .a (net558),
    .b (net561),
    .out (net656)
  );
  and_cell and133 (
    .a (net656),
    .b (net654),
    .out (net530)
  );
  and_cell and135 (
    .a (net655),
    .b (net654),
    .out (net636)
  );
  and_cell and136 (
    .a (net620),
    .b (net481),
    .out (net637)
  );
  and_cell and137 (
    .a (net621),
    .b (net481),
    .out (net639)
  );
  and_cell and138 (
    .a (net622),
    .b (net481),
    .out (net641)
  );
  and_cell and139 (
    .a (net623),
    .b (net481),
    .out (net643)
  );
  and_cell and140 (
    .a (net624),
    .b (net481),
    .out (net645)
  );
  and_cell and141 (
    .a (net625),
    .b (net481),
    .out (net647)
  );
  and_cell and142 (
    .a (net626),
    .b (net481),
    .out (net649)
  );
  and_cell and143 (
    .a (net627),
    .b (net481),
    .out (net651)
  );
  dffsr_cell flop84 (
    .d (net661),
    .clk (net1),
    .s (net662),
    .r (net104),
    .q (net26),
    .notq (net663)
  );
  mux_cell mux194 (
    .a (net26),
    .b (net664),
    .sel (net665),
    .out (net661)
  );
  xor_cell xor26 (
    .a (net101),
    .b (net481),
    .out (net667)
  );
  dffsr_cell flop85 (
    .d (net668),
    .clk (net1),
    .s (net669),
    .r (net104),
    .q (net28),
    .notq ()
  );
  mux_cell mux195 (
    .a (net670),
    .b (net28),
    .sel (net152),
    .out (net668)
  );
  not_cell not40 (
    .in (net671),
    .out (net670)
  );
  or_cell or55 (
    .a (net162),
    .b (net161),
    .out (net672)
  );
  or_cell or56 (
    .a (net160),
    .b (net159),
    .out (net673)
  );
  or_cell or57 (
    .a (net158),
    .b (net157),
    .out (net674)
  );
  or_cell or58 (
    .a (net156),
    .b (net151),
    .out (net675)
  );
  or_cell or59 (
    .a (net672),
    .b (net673),
    .out (net676)
  );
  or_cell or60 (
    .a (net674),
    .b (net675),
    .out (net677)
  );
  or_cell or61 (
    .a (net676),
    .b (net677),
    .out (net671)
  );
  xor_cell xor27 (
    .a (net678),
    .b (net122),
    .out (net120)
  );
  and_cell and144 (
    .a (net678),
    .b (net122),
    .out (net679)
  );
  xor_cell xor28 (
    .a (net125),
    .b (net679),
    .out (net124)
  );
  and_cell and145 (
    .a (net125),
    .b (net679),
    .out (net680)
  );
  xor_cell xor29 (
    .a (net128),
    .b (net680),
    .out (net127)
  );
  and_cell and146 (
    .a (net128),
    .b (net680),
    .out (net681)
  );
  xor_cell xor30 (
    .a (net131),
    .b (net681),
    .out (net130)
  );
  and_cell and147 (
    .a (net131),
    .b (net681),
    .out (net682)
  );
  xor_cell xor31 (
    .a (net134),
    .b (net682),
    .out (net133)
  );
  and_cell and148 (
    .a (net134),
    .b (net682),
    .out (net683)
  );
  xor_cell xor32 (
    .a (net137),
    .b (net683),
    .out (net136)
  );
  and_cell and149 (
    .a (net137),
    .b (net683),
    .out (net684)
  );
  xor_cell xor33 (
    .a (net140),
    .b (net684),
    .out (net139)
  );
  and_cell and150 (
    .a (net140),
    .b (net684),
    .out (net685)
  );
  xor_cell xor34 (
    .a (net143),
    .b (net685),
    .out (net142)
  );
  and_cell and151 (
    .a (net566),
    .b (net555),
    .out (net117)
  );
  and_cell and152 (
    .a (net555),
    .b (net400),
    .out (net686)
  );
  or_cell or62 (
    .a (net687),
    .b (net565),
    .out (net572)
  );
  and_cell and153 (
    .a (net656),
    .b (net686),
    .out (net688)
  );
  and_cell and154 (
    .a (net566),
    .b (net553),
    .out (net689)
  );
  nand_cell nand6 (
    .a (net689),
    .b (net688),
    .out (net690)
  );
  mux_cell mux197 (
    .a (net691),
    .b (net667),
    .sel (net690),
    .out (net692)
  );
  and_cell and157 (
    .a (net481),
    .b (net663),
    .out (net691)
  );
  mux_cell mux196 (
    .a (net692),
    .b (net693),
    .sel (net484),
    .out (net664)
  );
  mux_cell mux198 (
    .a (net94),
    .b (net35),
    .sel (net694),
    .out (net693)
  );
  mux_cell mux199 (
    .a (net38),
    .b (net695),
    .sel (net481),
    .out (net696)
  );
  mux_cell mux200 (
    .a (net49),
    .b (net35),
    .sel (net481),
    .out (net697)
  );
  mux_cell mux201 (
    .a (net58),
    .b (net38),
    .sel (net481),
    .out (net698)
  );
  mux_cell mux202 (
    .a (net67),
    .b (net49),
    .sel (net481),
    .out (net699)
  );
  mux_cell mux203 (
    .a (net76),
    .b (net58),
    .sel (net481),
    .out (net700)
  );
  mux_cell mux204 (
    .a (net85),
    .b (net67),
    .sel (net481),
    .out (net701)
  );
  mux_cell mux205 (
    .a (net94),
    .b (net76),
    .sel (net481),
    .out (net702)
  );
  mux_cell mux206 (
    .a (net703),
    .b (net85),
    .sel (net481),
    .out (net704)
  );
  mux_cell mux208 (
    .a (net705),
    .b (net26),
    .sel (net553),
    .out (net695)
  );
  mux_cell mux209 (
    .a (net706),
    .b (net26),
    .sel (net553),
    .out (net703)
  );
  and_cell and158 (
    .a (net484),
    .b (net94),
    .out (net706)
  );
  mux_cell mux207 (
    .a (net696),
    .b (net638),
    .sel (net556),
    .out (net529)
  );
  mux_cell mux210 (
    .a (net697),
    .b (net640),
    .sel (net556),
    .out (net532)
  );
  mux_cell mux211 (
    .a (net698),
    .b (net642),
    .sel (net556),
    .out (net534)
  );
  mux_cell mux212 (
    .a (net699),
    .b (net644),
    .sel (net556),
    .out (net536)
  );
  mux_cell mux213 (
    .a (net700),
    .b (net646),
    .sel (net556),
    .out (net538)
  );
  mux_cell mux214 (
    .a (net701),
    .b (net648),
    .sel (net556),
    .out (net540)
  );
  mux_cell mux215 (
    .a (net702),
    .b (net650),
    .sel (net556),
    .out (net542)
  );
  mux_cell mux216 (
    .a (net704),
    .b (net652),
    .sel (net556),
    .out (net544)
  );
  and_cell and134 (
    .a (net550),
    .b (net553),
    .out (net707)
  );
  and_cell and159 (
    .a (net688),
    .b (net707),
    .out (net687)
  );
  not_cell not41 (
    .in (net481),
    .out (net694)
  );
  and_cell and155 (
    .a (net711),
    .b (net712),
    .out (net665)
  );
  not_cell not42 (
    .in (net155),
    .out (net712)
  );
  or_cell or64 (
    .a (net713),
    .b (net714),
    .out (net715)
  );
  not_cell not43 (
    .in (net690),
    .out (net714)
  );
  or_cell or63 (
    .a (net715),
    .b (net563),
    .out (net711)
  );
  and_cell and156 (
    .a (net548),
    .b (net484),
    .out (net716)
  );
  and_cell and160 (
    .a (net552),
    .b (net566),
    .out (net717)
  );
  and_cell and161 (
    .a (net717),
    .b (net716),
    .out (net718)
  );
  and_cell and162 (
    .a (net718),
    .b (net688),
    .out (net713)
  );
endmodule
