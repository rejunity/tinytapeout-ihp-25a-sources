/*
 * Copyright (c) 2024 Sebastian Pfeiler
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_Qwendu_spi_fpu (
	  input  wire [7:0] ui_in,    // Dedicated inputs
	  output wire [7:0] uo_out,   // Dedicated outputs
	  input  wire [7:0] uio_in,   // IOs: Input path
	  output wire [7:0] uio_out,  // IOs: Output path
	  output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
	  input  wire       ena,      // always 1 when the design is powered, so you can ignore it
	  input  wire       clk,      // clock
	  input  wire       rst_n     // reset_n - low to reset
);
	assign uo_out[7:1]  = 7'b0;
	assign uio_out = 0;
	assign uio_oe  = 0;

	spi_fpu main(
		.clock(clk),
		.reset(!rst_n),
		.SPI_clock(ui_in[0]),
		.SPI_not_chip_select(ui_in[1]),
		.SPI_in(ui_in[2]),
		.SPI_out(uo_out[0])
	);
endmodule
