/* Automatically generated from https://wokwi.com/projects/414122607025630209 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_414122607025630209(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = ui_in[6];
  wire net3 = ui_in[7];
  wire net4;
  wire net5 = 1'b0;
  wire net6 = 1'b1;
  wire net7 = 1'b1;
  wire net8;
  wire net9;
  wire net10 = 1'b1;
  wire net11;
  wire net12;
  wire net13 = 1'b1;
  wire net14;
  wire net15;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19 = 1'b1;
  wire net20;
  wire net21;
  wire net22 = 1'b0;
  wire net23;
  wire net24;
  wire net25 = 1'b1;
  wire net26;
  wire net27;
  wire net28 = 1'b1;
  wire net29;
  wire net30;
  wire net31 = 1'b0;
  wire net32;
  wire net33;
  wire net34 = 1'b0;
  wire net35;
  wire net36;
  wire net37 = 1'b1;
  wire net38;
  wire net39;
  wire net40 = 1'b0;
  wire net41;
  wire net42;
  wire net43 = 1'b1;
  wire net44;
  wire net45;
  wire net46 = 1'b0;
  wire net47;
  wire net48;
  wire net49 = 1'b1;
  wire net50;
  wire net51;
  wire net52 = 1'b1;
  wire net53;
  wire net54;
  wire net55 = 1'b1;
  wire net56;
  wire net57;
  wire net58 = 1'b1;
  wire net59;
  wire net60 = 1'b0;
  wire net61 = 1'b0;
  wire net62 = 1'b0;
  wire net63;
  wire net64;
  wire net65 = 1'b1;
  wire net66;
  wire net67;
  wire net68 = 1'b1;
  wire net69;
  wire net70;
  wire net71 = 1'b1;
  wire net72;
  wire net73;
  wire net74 = 1'b1;
  wire net75;
  wire net76;
  wire net77 = 1'b0;
  wire net78;
  wire net79;
  wire net80 = 1'b0;
  wire net81;
  wire net82;
  wire net83 = 1'b0;
  wire net84;
  wire net85;
  wire net86 = 1'b0;
  wire net87;
  wire net88;
  wire net89 = 1'b1;
  wire net90;
  wire net91;
  wire net92 = 1'b0;
  wire net93;
  wire net94;
  wire net95 = 1'b0;
  wire net96;
  wire net97;
  wire net98 = 1'b1;
  wire net99;
  wire net100;
  wire net101 = 1'b0;
  wire net102;
  wire net103;
  wire net104 = 1'b1;
  wire net105;
  wire net106;
  wire net107 = 1'b1;
  wire net108;
  wire net109;
  wire net110 = 1'b1;
  wire net111;
  wire net112;
  wire net113 = 1'b1;
  wire net114;
  wire net115 = 1'b0;
  wire net116;
  wire net117 = 1'b1;
  wire net118;
  wire net119;
  wire net120 = 1'b1;
  wire net121;
  wire net122;
  wire net123 = 1'b1;
  wire net124;
  wire net125;
  wire net126 = 1'b1;
  wire net127;
  wire net128;
  wire net129 = 1'b1;
  wire net130;
  wire net131;
  wire net132 = 1'b1;
  wire net133;
  wire net134;
  wire net135 = 1'b1;
  wire net136;
  wire net137;
  wire net138 = 1'b1;
  wire net139;
  wire net140;
  wire net141 = 1'b1;
  wire net142;
  wire net143;
  wire net144 = 1'b1;
  wire net145;
  wire net146;
  wire net147 = 1'b1;
  wire net148;
  wire net149;
  wire net150 = 1'b1;
  wire net151;
  wire net152;
  wire net153 = 1'b0;
  wire net154;
  wire net155;
  wire net156 = 1'b1;
  wire net157;
  wire net158;
  wire net159 = 1'b0;
  wire net160;
  wire net161;
  wire net162 = 1'b0;
  wire net163;
  wire net164;
  wire net165 = 1'b0;
  wire net166;
  wire net167;
  wire net168 = 1'b0;
  wire net169;
  wire net170;
  wire net171 = 1'b0;
  wire net172;
  wire net173;
  wire net174 = 1'b1;
  wire net175;
  wire net176;
  wire net177 = 1'b0;
  wire net178;
  wire net179;
  wire net180 = 1'b1;
  wire net181;
  wire net182;
  wire net183 = 1'b1;
  wire net184;
  wire net185;
  wire net186 = 1'b1;
  wire net187;
  wire net188;
  wire net189 = 1'b1;
  wire net190;
  wire net191 = 1'b0;
  wire net192;
  wire net193 = 1'b1;
  wire net194;
  wire net195;
  wire net196 = 1'b1;
  wire net197;
  wire net198;
  wire net199 = 1'b1;
  wire net200;
  wire net201;
  wire net202 = 1'b1;
  wire net203;
  wire net204;
  wire net205 = 1'b1;
  wire net206;
  wire net207;
  wire net208 = 1'b1;
  wire net209;
  wire net210;
  wire net211 = 1'b1;
  wire net212;
  wire net213;
  wire net214 = 1'b1;
  wire net215;
  wire net216;
  wire net217 = 1'b0;
  wire net218;
  wire net219;
  wire net220 = 1'b1;
  wire net221;
  wire net222;
  wire net223 = 1'b1;
  wire net224;
  wire net225;
  wire net226 = 1'b1;
  wire net227;
  wire net228;
  wire net229 = 1'b1;
  wire net230;
  wire net231;
  wire net232 = 1'b0;
  wire net233;
  wire net234;
  wire net235 = 1'b0;
  wire net236;
  wire net237;
  wire net238 = 1'b1;
  wire net239;
  wire net240;
  wire net241 = 1'b0;
  wire net242;
  wire net243;
  wire net244 = 1'b1;
  wire net245;
  wire net246;
  wire net247 = 1'b1;
  wire net248;
  wire net249;
  wire net250 = 1'b1;
  wire net251;
  wire net252;
  wire net253 = 1'b1;
  wire net254;
  wire net255 = 1'b0;
  wire net256;
  wire net257 = 1'b1;
  wire net258;
  wire net259;
  wire net260 = 1'b1;
  wire net261;
  wire net262;
  wire net263 = 1'b1;
  wire net264;
  wire net265;
  wire net266 = 1'b1;
  wire net267;
  wire net268;
  wire net269 = 1'b1;
  wire net270;
  wire net271;
  wire net272 = 1'b1;
  wire net273;
  wire net274;
  wire net275 = 1'b1;
  wire net276;
  wire net277;
  wire net278 = 1'b1;
  wire net279;
  wire net280;
  wire net281 = 1'b0;
  wire net282;
  wire net283;
  wire net284 = 1'b1;
  wire net285;
  wire net286;
  wire net287 = 1'b1;
  wire net288;
  wire net289;
  wire net290 = 1'b0;
  wire net291;
  wire net292;
  wire net293 = 1'b1;
  wire net294;
  wire net295;
  wire net296 = 1'b0;
  wire net297;
  wire net298;
  wire net299 = 1'b0;
  wire net300;
  wire net301;
  wire net302 = 1'b1;
  wire net303;
  wire net304;
  wire net305 = 1'b0;
  wire net306;
  wire net307;
  wire net308 = 1'b1;
  wire net309;
  wire net310;
  wire net311 = 1'b1;
  wire net312;
  wire net313;
  wire net314 = 1'b1;
  wire net315;
  wire net316;
  wire net317 = 1'b1;
  wire net318;
  wire net319 = 1'b0;
  wire net320;
  wire net321 = 1'b1;
  wire net322;
  wire net323;
  wire net324 = 1'b1;
  wire net325;
  wire net326;
  wire net327 = 1'b1;
  wire net328;
  wire net329;
  wire net330 = 1'b1;
  wire net331 = 1'b1;
  wire net332;
  wire net333;
  wire net334 = 1'b1;
  wire net335;
  wire net336;
  wire net337 = 1'b1;
  wire net338;
  wire net339;
  wire net340 = 1'b1;
  wire net341;
  wire net342;
  wire net343 = 1'b1;
  wire net344;
  wire net345;
  wire net346 = 1'b0;
  wire net347;
  wire net348;
  wire net349 = 1'b1;
  wire net350;
  wire net351;
  wire net352 = 1'b0;
  wire net353;
  wire net354;
  wire net355 = 1'b0;
  wire net356;
  wire net357;
  wire net358 = 1'b0;
  wire net359;
  wire net360;
  wire net361 = 1'b0;
  wire net362;
  wire net363;
  wire net364 = 1'b0;
  wire net365;
  wire net366;
  wire net367 = 1'b1;
  wire net368;
  wire net369;
  wire net370 = 1'b0;
  wire net371;
  wire net372;
  wire net373 = 1'b1;
  wire net374;
  wire net375;
  wire net376 = 1'b1;
  wire net377;
  wire net378;
  wire net379 = 1'b1;
  wire net380;
  wire net381;
  wire net382 = 1'b1;
  wire net383;
  wire net384 = 1'b0;
  wire net385;
  wire net386 = 1'b1;
  wire net387;
  wire net388;
  wire net389 = 1'b1;
  wire net390;
  wire net391;
  wire net392 = 1'b1;
  wire net393;
  wire net394;
  wire net395 = 1'b1;
  wire net396;
  wire net397;
  wire net398 = 1'b1;
  wire net399;
  wire net400;
  wire net401 = 1'b1;
  wire net402;
  wire net403;
  wire net404 = 1'b1;
  wire net405;
  wire net406;
  wire net407 = 1'b1;
  wire net408;
  wire net409;
  wire net410 = 1'b0;
  wire net411;
  wire net412;
  wire net413 = 1'b1;
  wire net414;
  wire net415;
  wire net416 = 1'b0;
  wire net417;
  wire net418;
  wire net419 = 1'b0;
  wire net420;
  wire net421;
  wire net422 = 1'b1;
  wire net423;
  wire net424;
  wire net425 = 1'b0;
  wire net426;
  wire net427;
  wire net428 = 1'b0;
  wire net429;
  wire net430;
  wire net431 = 1'b1;
  wire net432;
  wire net433;
  wire net434 = 1'b0;
  wire net435;
  wire net436;
  wire net437 = 1'b1;
  wire net438;
  wire net439;
  wire net440 = 1'b1;
  wire net441;
  wire net442;
  wire net443 = 1'b1;
  wire net444;
  wire net445;
  wire net446 = 1'b1;
  wire net447;
  wire net448 = 1'b0;
  wire net449;
  wire net450 = 1'b1;
  wire net451;
  wire net452;
  wire net453 = 1'b1;
  wire net454;
  wire net455;
  wire net456 = 1'b1;
  wire net457;
  wire net458;
  wire net459 = 1'b1;
  wire net460;
  wire net461;
  wire net462 = 1'b1;
  wire net463;
  wire net464;
  wire net465 = 1'b1;
  wire net466;
  wire net467;
  wire net468 = 1'b1;
  wire net469;
  wire net470;
  wire net471 = 1'b1;
  wire net472;
  wire net473;
  wire net474 = 1'b0;
  wire net475;
  wire net476;
  wire net477 = 1'b0;
  wire net478;
  wire net479;
  wire net480 = 1'b1;
  wire net481;
  wire net482;
  wire net483 = 1'b0;
  wire net484;
  wire net485;
  wire net486 = 1'b1;
  wire net487;
  wire net488;
  wire net489 = 1'b0;
  wire net490;
  wire net491;
  wire net492 = 1'b0;
  wire net493;
  wire net494;
  wire net495 = 1'b0;
  wire net496;
  wire net497;
  wire net498 = 1'b0;
  wire net499;
  wire net500;
  wire net501 = 1'b1;
  wire net502;
  wire net503;
  wire net504 = 1'b1;
  wire net505;
  wire net506;
  wire net507 = 1'b1;
  wire net508;
  wire net509;
  wire net510 = 1'b1;
  wire net511 = 1'b0;
  wire net512;
  wire net513 = 1'b1;
  wire net514;
  wire net515;
  wire net516 = 1'b1;
  wire net517;
  wire net518;
  wire net519 = 1'b1;
  wire net520;
  wire net521;
  wire net522 = 1'b1;

  assign uo_out[0] = net3;
  assign uo_out[1] = net2;
  assign uo_out[2] = 0;
  assign uo_out[3] = 0;
  assign uo_out[4] = 0;
  assign uo_out[5] = 0;
  assign uo_out[6] = 0;
  assign uo_out[7] = net4;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  dff_cell flop1 (
    .d (net8),
    .clk (net1),
    .q (net9),
    .notq ()
  );
  mux_cell mux1 (
    .a (net10),
    .b (net11),
    .sel (net2),
    .out (net8)
  );
  dff_cell flop3 (
    .d (net12),
    .clk (net1),
    .q (net11),
    .notq ()
  );
  mux_cell mux3 (
    .a (net13),
    .b (net14),
    .sel (net2),
    .out (net12)
  );
  dff_cell flop4 (
    .d (net15),
    .clk (net1),
    .q (net14),
    .notq ()
  );
  mux_cell mux4 (
    .a (net16),
    .b (net17),
    .sel (net2),
    .out (net15)
  );
  dff_cell flop5 (
    .d (net18),
    .clk (net1),
    .q (net17),
    .notq ()
  );
  mux_cell mux5 (
    .a (net19),
    .b (net20),
    .sel (net2),
    .out (net18)
  );
  dff_cell flop6 (
    .d (net21),
    .clk (net1),
    .q (net20),
    .notq ()
  );
  mux_cell mux6 (
    .a (net22),
    .b (net23),
    .sel (net2),
    .out (net21)
  );
  dff_cell flop7 (
    .d (net24),
    .clk (net1),
    .q (net23),
    .notq ()
  );
  mux_cell mux7 (
    .a (net25),
    .b (net26),
    .sel (net2),
    .out (net24)
  );
  dff_cell flop8 (
    .d (net27),
    .clk (net1),
    .q (net26),
    .notq ()
  );
  mux_cell mux8 (
    .a (net28),
    .b (net29),
    .sel (net2),
    .out (net27)
  );
  dff_cell flop9 (
    .d (net30),
    .clk (net1),
    .q (net29),
    .notq ()
  );
  mux_cell mux9 (
    .a (net31),
    .b (net32),
    .sel (net2),
    .out (net30)
  );
  dff_cell flop10 (
    .d (net33),
    .clk (net1),
    .q (net32),
    .notq ()
  );
  mux_cell mux10 (
    .a (net34),
    .b (net35),
    .sel (net2),
    .out (net33)
  );
  dff_cell flop11 (
    .d (net36),
    .clk (net1),
    .q (net35),
    .notq ()
  );
  mux_cell mux11 (
    .a (net37),
    .b (net38),
    .sel (net2),
    .out (net36)
  );
  dff_cell flop12 (
    .d (net39),
    .clk (net1),
    .q (net38),
    .notq ()
  );
  mux_cell mux12 (
    .a (net40),
    .b (net41),
    .sel (net2),
    .out (net39)
  );
  dff_cell flop13 (
    .d (net42),
    .clk (net1),
    .q (net41),
    .notq ()
  );
  mux_cell mux13 (
    .a (net43),
    .b (net44),
    .sel (net2),
    .out (net42)
  );
  dff_cell flop14 (
    .d (net45),
    .clk (net1),
    .q (net44),
    .notq ()
  );
  mux_cell mux14 (
    .a (net46),
    .b (net47),
    .sel (net2),
    .out (net45)
  );
  dff_cell flop15 (
    .d (net48),
    .clk (net1),
    .q (net47),
    .notq ()
  );
  mux_cell mux15 (
    .a (net49),
    .b (net50),
    .sel (net2),
    .out (net48)
  );
  dff_cell flop16 (
    .d (net51),
    .clk (net1),
    .q (net50),
    .notq ()
  );
  mux_cell mux16 (
    .a (net52),
    .b (net53),
    .sel (net2),
    .out (net51)
  );
  dff_cell flop17 (
    .d (net54),
    .clk (net1),
    .q (net53),
    .notq ()
  );
  mux_cell mux17 (
    .a (net55),
    .b (net56),
    .sel (net2),
    .out (net54)
  );
  dff_cell flop18 (
    .d (net57),
    .clk (net1),
    .q (net56),
    .notq ()
  );
  mux_cell mux18 (
    .a (net58),
    .b (net59),
    .sel (net2),
    .out (net57)
  );
  dff_cell flop2 (
    .d (net63),
    .clk (net1),
    .q (net64),
    .notq ()
  );
  mux_cell mux19 (
    .a (net65),
    .b (net66),
    .sel (net2),
    .out (net63)
  );
  dff_cell flop19 (
    .d (net67),
    .clk (net1),
    .q (net66),
    .notq ()
  );
  mux_cell mux20 (
    .a (net68),
    .b (net69),
    .sel (net2),
    .out (net67)
  );
  dff_cell flop20 (
    .d (net70),
    .clk (net1),
    .q (net69),
    .notq ()
  );
  mux_cell mux21 (
    .a (net71),
    .b (net72),
    .sel (net2),
    .out (net70)
  );
  dff_cell flop21 (
    .d (net73),
    .clk (net1),
    .q (net72),
    .notq ()
  );
  mux_cell mux22 (
    .a (net74),
    .b (net75),
    .sel (net2),
    .out (net73)
  );
  dff_cell flop22 (
    .d (net76),
    .clk (net1),
    .q (net75),
    .notq ()
  );
  mux_cell mux23 (
    .a (net77),
    .b (net78),
    .sel (net2),
    .out (net76)
  );
  dff_cell flop23 (
    .d (net79),
    .clk (net1),
    .q (net78),
    .notq ()
  );
  mux_cell mux24 (
    .a (net80),
    .b (net81),
    .sel (net2),
    .out (net79)
  );
  dff_cell flop24 (
    .d (net82),
    .clk (net1),
    .q (net81),
    .notq ()
  );
  mux_cell mux25 (
    .a (net83),
    .b (net84),
    .sel (net2),
    .out (net82)
  );
  dff_cell flop25 (
    .d (net85),
    .clk (net1),
    .q (net84),
    .notq ()
  );
  mux_cell mux26 (
    .a (net86),
    .b (net87),
    .sel (net2),
    .out (net85)
  );
  dff_cell flop26 (
    .d (net88),
    .clk (net1),
    .q (net87),
    .notq ()
  );
  mux_cell mux27 (
    .a (net89),
    .b (net90),
    .sel (net2),
    .out (net88)
  );
  dff_cell flop27 (
    .d (net91),
    .clk (net1),
    .q (net90),
    .notq ()
  );
  mux_cell mux28 (
    .a (net92),
    .b (net93),
    .sel (net2),
    .out (net91)
  );
  dff_cell flop28 (
    .d (net94),
    .clk (net1),
    .q (net93),
    .notq ()
  );
  mux_cell mux29 (
    .a (net95),
    .b (net96),
    .sel (net2),
    .out (net94)
  );
  dff_cell flop29 (
    .d (net97),
    .clk (net1),
    .q (net96),
    .notq ()
  );
  mux_cell mux30 (
    .a (net98),
    .b (net99),
    .sel (net2),
    .out (net97)
  );
  dff_cell flop30 (
    .d (net100),
    .clk (net1),
    .q (net99),
    .notq ()
  );
  mux_cell mux31 (
    .a (net101),
    .b (net102),
    .sel (net2),
    .out (net100)
  );
  dff_cell flop31 (
    .d (net103),
    .clk (net1),
    .q (net102),
    .notq ()
  );
  mux_cell mux32 (
    .a (net104),
    .b (net105),
    .sel (net2),
    .out (net103)
  );
  dff_cell flop32 (
    .d (net106),
    .clk (net1),
    .q (net105),
    .notq ()
  );
  mux_cell mux33 (
    .a (net107),
    .b (net108),
    .sel (net2),
    .out (net106)
  );
  dff_cell flop33 (
    .d (net109),
    .clk (net1),
    .q (net108),
    .notq ()
  );
  mux_cell mux34 (
    .a (net110),
    .b (net111),
    .sel (net2),
    .out (net109)
  );
  dff_cell flop34 (
    .d (net112),
    .clk (net1),
    .q (net111),
    .notq ()
  );
  mux_cell mux35 (
    .a (net113),
    .b (net114),
    .sel (net2),
    .out (net112)
  );
  dff_cell flop35 (
    .d (net116),
    .clk (net1),
    .q (net59),
    .notq ()
  );
  mux_cell mux36 (
    .a (net117),
    .b (net118),
    .sel (net2),
    .out (net116)
  );
  dff_cell flop36 (
    .d (net119),
    .clk (net1),
    .q (net118),
    .notq ()
  );
  mux_cell mux37 (
    .a (net120),
    .b (net121),
    .sel (net2),
    .out (net119)
  );
  dff_cell flop37 (
    .d (net122),
    .clk (net1),
    .q (net121),
    .notq ()
  );
  mux_cell mux38 (
    .a (net123),
    .b (net124),
    .sel (net2),
    .out (net122)
  );
  dff_cell flop38 (
    .d (net125),
    .clk (net1),
    .q (net124),
    .notq ()
  );
  mux_cell mux39 (
    .a (net126),
    .b (net64),
    .sel (net2),
    .out (net125)
  );
  dff_cell flop39 (
    .d (net127),
    .clk (net1),
    .q (net128),
    .notq ()
  );
  mux_cell mux40 (
    .a (net129),
    .b (net130),
    .sel (net2),
    .out (net127)
  );
  dff_cell flop40 (
    .d (net131),
    .clk (net1),
    .q (net130),
    .notq ()
  );
  mux_cell mux41 (
    .a (net132),
    .b (net133),
    .sel (net2),
    .out (net131)
  );
  dff_cell flop41 (
    .d (net134),
    .clk (net1),
    .q (net133),
    .notq ()
  );
  mux_cell mux42 (
    .a (net135),
    .b (net136),
    .sel (net2),
    .out (net134)
  );
  dff_cell flop42 (
    .d (net137),
    .clk (net1),
    .q (net136),
    .notq ()
  );
  mux_cell mux43 (
    .a (net138),
    .b (net9),
    .sel (net2),
    .out (net137)
  );
  dff_cell flop43 (
    .d (net139),
    .clk (net1),
    .q (net140),
    .notq ()
  );
  mux_cell mux44 (
    .a (net141),
    .b (net142),
    .sel (net2),
    .out (net139)
  );
  dff_cell flop44 (
    .d (net143),
    .clk (net1),
    .q (net142),
    .notq ()
  );
  mux_cell mux45 (
    .a (net144),
    .b (net145),
    .sel (net2),
    .out (net143)
  );
  dff_cell flop45 (
    .d (net146),
    .clk (net1),
    .q (net145),
    .notq ()
  );
  mux_cell mux46 (
    .a (net147),
    .b (net148),
    .sel (net2),
    .out (net146)
  );
  dff_cell flop46 (
    .d (net149),
    .clk (net1),
    .q (net148),
    .notq ()
  );
  mux_cell mux47 (
    .a (net150),
    .b (net151),
    .sel (net2),
    .out (net149)
  );
  dff_cell flop47 (
    .d (net152),
    .clk (net1),
    .q (net151),
    .notq ()
  );
  mux_cell mux48 (
    .a (net153),
    .b (net154),
    .sel (net2),
    .out (net152)
  );
  dff_cell flop48 (
    .d (net155),
    .clk (net1),
    .q (net154),
    .notq ()
  );
  mux_cell mux49 (
    .a (net156),
    .b (net157),
    .sel (net2),
    .out (net155)
  );
  dff_cell flop49 (
    .d (net158),
    .clk (net1),
    .q (net157),
    .notq ()
  );
  mux_cell mux50 (
    .a (net159),
    .b (net160),
    .sel (net2),
    .out (net158)
  );
  dff_cell flop50 (
    .d (net161),
    .clk (net1),
    .q (net160),
    .notq ()
  );
  mux_cell mux51 (
    .a (net162),
    .b (net163),
    .sel (net2),
    .out (net161)
  );
  dff_cell flop51 (
    .d (net164),
    .clk (net1),
    .q (net163),
    .notq ()
  );
  mux_cell mux52 (
    .a (net165),
    .b (net166),
    .sel (net2),
    .out (net164)
  );
  dff_cell flop52 (
    .d (net167),
    .clk (net1),
    .q (net166),
    .notq ()
  );
  mux_cell mux53 (
    .a (net168),
    .b (net169),
    .sel (net2),
    .out (net167)
  );
  dff_cell flop53 (
    .d (net170),
    .clk (net1),
    .q (net169),
    .notq ()
  );
  mux_cell mux54 (
    .a (net171),
    .b (net172),
    .sel (net2),
    .out (net170)
  );
  dff_cell flop54 (
    .d (net173),
    .clk (net1),
    .q (net172),
    .notq ()
  );
  mux_cell mux55 (
    .a (net174),
    .b (net175),
    .sel (net2),
    .out (net173)
  );
  dff_cell flop55 (
    .d (net176),
    .clk (net1),
    .q (net175),
    .notq ()
  );
  mux_cell mux56 (
    .a (net177),
    .b (net178),
    .sel (net2),
    .out (net176)
  );
  dff_cell flop56 (
    .d (net179),
    .clk (net1),
    .q (net178),
    .notq ()
  );
  mux_cell mux57 (
    .a (net180),
    .b (net181),
    .sel (net2),
    .out (net179)
  );
  dff_cell flop57 (
    .d (net182),
    .clk (net1),
    .q (net181),
    .notq ()
  );
  mux_cell mux58 (
    .a (net183),
    .b (net184),
    .sel (net2),
    .out (net182)
  );
  dff_cell flop58 (
    .d (net185),
    .clk (net1),
    .q (net184),
    .notq ()
  );
  mux_cell mux59 (
    .a (net186),
    .b (net187),
    .sel (net2),
    .out (net185)
  );
  dff_cell flop59 (
    .d (net188),
    .clk (net1),
    .q (net187),
    .notq ()
  );
  mux_cell mux60 (
    .a (net189),
    .b (net190),
    .sel (net2),
    .out (net188)
  );
  dff_cell flop60 (
    .d (net192),
    .clk (net1),
    .q (net114),
    .notq ()
  );
  mux_cell mux61 (
    .a (net193),
    .b (net194),
    .sel (net2),
    .out (net192)
  );
  dff_cell flop61 (
    .d (net195),
    .clk (net1),
    .q (net194),
    .notq ()
  );
  mux_cell mux62 (
    .a (net196),
    .b (net197),
    .sel (net2),
    .out (net195)
  );
  dff_cell flop62 (
    .d (net198),
    .clk (net1),
    .q (net197),
    .notq ()
  );
  mux_cell mux63 (
    .a (net199),
    .b (net200),
    .sel (net2),
    .out (net198)
  );
  dff_cell flop63 (
    .d (net201),
    .clk (net1),
    .q (net200),
    .notq ()
  );
  mux_cell mux64 (
    .a (net202),
    .b (net140),
    .sel (net2),
    .out (net201)
  );
  dff_cell flop64 (
    .d (net203),
    .clk (net1),
    .q (net204),
    .notq ()
  );
  mux_cell mux65 (
    .a (net205),
    .b (net206),
    .sel (net2),
    .out (net203)
  );
  dff_cell flop65 (
    .d (net207),
    .clk (net1),
    .q (net206),
    .notq ()
  );
  mux_cell mux66 (
    .a (net208),
    .b (net209),
    .sel (net2),
    .out (net207)
  );
  dff_cell flop66 (
    .d (net210),
    .clk (net1),
    .q (net209),
    .notq ()
  );
  mux_cell mux67 (
    .a (net211),
    .b (net212),
    .sel (net2),
    .out (net210)
  );
  dff_cell flop67 (
    .d (net213),
    .clk (net1),
    .q (net212),
    .notq ()
  );
  mux_cell mux68 (
    .a (net214),
    .b (net215),
    .sel (net2),
    .out (net213)
  );
  dff_cell flop68 (
    .d (net216),
    .clk (net1),
    .q (net215),
    .notq ()
  );
  mux_cell mux69 (
    .a (net217),
    .b (net218),
    .sel (net2),
    .out (net216)
  );
  dff_cell flop69 (
    .d (net219),
    .clk (net1),
    .q (net218),
    .notq ()
  );
  mux_cell mux70 (
    .a (net220),
    .b (net221),
    .sel (net2),
    .out (net219)
  );
  dff_cell flop70 (
    .d (net222),
    .clk (net1),
    .q (net221),
    .notq ()
  );
  mux_cell mux71 (
    .a (net223),
    .b (net224),
    .sel (net2),
    .out (net222)
  );
  dff_cell flop71 (
    .d (net225),
    .clk (net1),
    .q (net224),
    .notq ()
  );
  mux_cell mux72 (
    .a (net226),
    .b (net227),
    .sel (net2),
    .out (net225)
  );
  dff_cell flop72 (
    .d (net228),
    .clk (net1),
    .q (net227),
    .notq ()
  );
  mux_cell mux73 (
    .a (net229),
    .b (net230),
    .sel (net2),
    .out (net228)
  );
  dff_cell flop73 (
    .d (net231),
    .clk (net1),
    .q (net230),
    .notq ()
  );
  mux_cell mux74 (
    .a (net232),
    .b (net233),
    .sel (net2),
    .out (net231)
  );
  dff_cell flop74 (
    .d (net234),
    .clk (net1),
    .q (net233),
    .notq ()
  );
  mux_cell mux75 (
    .a (net235),
    .b (net236),
    .sel (net2),
    .out (net234)
  );
  dff_cell flop75 (
    .d (net237),
    .clk (net1),
    .q (net236),
    .notq ()
  );
  mux_cell mux76 (
    .a (net238),
    .b (net239),
    .sel (net2),
    .out (net237)
  );
  dff_cell flop76 (
    .d (net240),
    .clk (net1),
    .q (net239),
    .notq ()
  );
  mux_cell mux77 (
    .a (net241),
    .b (net242),
    .sel (net2),
    .out (net240)
  );
  dff_cell flop77 (
    .d (net243),
    .clk (net1),
    .q (net242),
    .notq ()
  );
  mux_cell mux78 (
    .a (net244),
    .b (net245),
    .sel (net2),
    .out (net243)
  );
  dff_cell flop78 (
    .d (net246),
    .clk (net1),
    .q (net245),
    .notq ()
  );
  mux_cell mux79 (
    .a (net247),
    .b (net248),
    .sel (net2),
    .out (net246)
  );
  dff_cell flop79 (
    .d (net249),
    .clk (net1),
    .q (net248),
    .notq ()
  );
  mux_cell mux80 (
    .a (net250),
    .b (net251),
    .sel (net2),
    .out (net249)
  );
  dff_cell flop80 (
    .d (net252),
    .clk (net1),
    .q (net251),
    .notq ()
  );
  mux_cell mux81 (
    .a (net253),
    .b (net254),
    .sel (net2),
    .out (net252)
  );
  dff_cell flop81 (
    .d (net256),
    .clk (net1),
    .q (net190),
    .notq ()
  );
  mux_cell mux82 (
    .a (net257),
    .b (net258),
    .sel (net2),
    .out (net256)
  );
  dff_cell flop82 (
    .d (net259),
    .clk (net1),
    .q (net258),
    .notq ()
  );
  mux_cell mux83 (
    .a (net260),
    .b (net261),
    .sel (net2),
    .out (net259)
  );
  dff_cell flop83 (
    .d (net262),
    .clk (net1),
    .q (net261),
    .notq ()
  );
  mux_cell mux84 (
    .a (net263),
    .b (net264),
    .sel (net2),
    .out (net262)
  );
  dff_cell flop84 (
    .d (net265),
    .clk (net1),
    .q (net264),
    .notq ()
  );
  mux_cell mux85 (
    .a (net266),
    .b (net204),
    .sel (net2),
    .out (net265)
  );
  dff_cell flop85 (
    .d (net267),
    .clk (net1),
    .q (net268),
    .notq ()
  );
  mux_cell mux86 (
    .a (net269),
    .b (net270),
    .sel (net2),
    .out (net267)
  );
  dff_cell flop86 (
    .d (net271),
    .clk (net1),
    .q (net270),
    .notq ()
  );
  mux_cell mux87 (
    .a (net272),
    .b (net273),
    .sel (net2),
    .out (net271)
  );
  dff_cell flop87 (
    .d (net274),
    .clk (net1),
    .q (net273),
    .notq ()
  );
  mux_cell mux88 (
    .a (net275),
    .b (net276),
    .sel (net2),
    .out (net274)
  );
  dff_cell flop88 (
    .d (net277),
    .clk (net1),
    .q (net276),
    .notq ()
  );
  mux_cell mux89 (
    .a (net278),
    .b (net279),
    .sel (net2),
    .out (net277)
  );
  dff_cell flop89 (
    .d (net280),
    .clk (net1),
    .q (net279),
    .notq ()
  );
  mux_cell mux90 (
    .a (net281),
    .b (net282),
    .sel (net2),
    .out (net280)
  );
  dff_cell flop90 (
    .d (net283),
    .clk (net1),
    .q (net282),
    .notq ()
  );
  mux_cell mux91 (
    .a (net284),
    .b (net285),
    .sel (net2),
    .out (net283)
  );
  dff_cell flop91 (
    .d (net286),
    .clk (net1),
    .q (net285),
    .notq ()
  );
  mux_cell mux92 (
    .a (net287),
    .b (net288),
    .sel (net2),
    .out (net286)
  );
  dff_cell flop92 (
    .d (net289),
    .clk (net1),
    .q (net288),
    .notq ()
  );
  mux_cell mux93 (
    .a (net290),
    .b (net291),
    .sel (net2),
    .out (net289)
  );
  dff_cell flop93 (
    .d (net292),
    .clk (net1),
    .q (net291),
    .notq ()
  );
  mux_cell mux94 (
    .a (net293),
    .b (net294),
    .sel (net2),
    .out (net292)
  );
  dff_cell flop94 (
    .d (net295),
    .clk (net1),
    .q (net294),
    .notq ()
  );
  mux_cell mux95 (
    .a (net296),
    .b (net297),
    .sel (net2),
    .out (net295)
  );
  dff_cell flop95 (
    .d (net298),
    .clk (net1),
    .q (net297),
    .notq ()
  );
  mux_cell mux96 (
    .a (net299),
    .b (net300),
    .sel (net2),
    .out (net298)
  );
  dff_cell flop96 (
    .d (net301),
    .clk (net1),
    .q (net300),
    .notq ()
  );
  mux_cell mux97 (
    .a (net302),
    .b (net303),
    .sel (net2),
    .out (net301)
  );
  dff_cell flop97 (
    .d (net304),
    .clk (net1),
    .q (net303),
    .notq ()
  );
  mux_cell mux98 (
    .a (net305),
    .b (net306),
    .sel (net2),
    .out (net304)
  );
  dff_cell flop98 (
    .d (net307),
    .clk (net1),
    .q (net306),
    .notq ()
  );
  mux_cell mux99 (
    .a (net308),
    .b (net309),
    .sel (net2),
    .out (net307)
  );
  dff_cell flop99 (
    .d (net310),
    .clk (net1),
    .q (net309),
    .notq ()
  );
  mux_cell mux100 (
    .a (net311),
    .b (net312),
    .sel (net2),
    .out (net310)
  );
  dff_cell flop100 (
    .d (net313),
    .clk (net1),
    .q (net312),
    .notq ()
  );
  mux_cell mux101 (
    .a (net314),
    .b (net315),
    .sel (net2),
    .out (net313)
  );
  dff_cell flop101 (
    .d (net316),
    .clk (net1),
    .q (net315),
    .notq ()
  );
  mux_cell mux102 (
    .a (net317),
    .b (net318),
    .sel (net2),
    .out (net316)
  );
  dff_cell flop102 (
    .d (net320),
    .clk (net1),
    .q (net254),
    .notq ()
  );
  mux_cell mux103 (
    .a (net321),
    .b (net322),
    .sel (net2),
    .out (net320)
  );
  dff_cell flop103 (
    .d (net323),
    .clk (net1),
    .q (net322),
    .notq ()
  );
  mux_cell mux104 (
    .a (net324),
    .b (net325),
    .sel (net2),
    .out (net323)
  );
  dff_cell flop104 (
    .d (net326),
    .clk (net1),
    .q (net325),
    .notq ()
  );
  mux_cell mux105 (
    .a (net327),
    .b (net328),
    .sel (net2),
    .out (net326)
  );
  dff_cell flop105 (
    .d (net329),
    .clk (net1),
    .q (net328),
    .notq ()
  );
  mux_cell mux106 (
    .a (net330),
    .b (net268),
    .sel (net2),
    .out (net329)
  );
  mux_cell mux2 (
    .a (net331),
    .b (net128),
    .sel (net3),
    .out (net4)
  );
  dff_cell flop106 (
    .d (net332),
    .clk (net1),
    .q (net333),
    .notq ()
  );
  mux_cell mux107 (
    .a (net334),
    .b (net335),
    .sel (net2),
    .out (net332)
  );
  dff_cell flop107 (
    .d (net336),
    .clk (net1),
    .q (net335),
    .notq ()
  );
  mux_cell mux108 (
    .a (net337),
    .b (net338),
    .sel (net2),
    .out (net336)
  );
  dff_cell flop108 (
    .d (net339),
    .clk (net1),
    .q (net338),
    .notq ()
  );
  mux_cell mux109 (
    .a (net340),
    .b (net341),
    .sel (net2),
    .out (net339)
  );
  dff_cell flop109 (
    .d (net342),
    .clk (net1),
    .q (net341),
    .notq ()
  );
  mux_cell mux110 (
    .a (net343),
    .b (net344),
    .sel (net2),
    .out (net342)
  );
  dff_cell flop110 (
    .d (net345),
    .clk (net1),
    .q (net344),
    .notq ()
  );
  mux_cell mux111 (
    .a (net346),
    .b (net347),
    .sel (net2),
    .out (net345)
  );
  dff_cell flop111 (
    .d (net348),
    .clk (net1),
    .q (net347),
    .notq ()
  );
  mux_cell mux112 (
    .a (net349),
    .b (net350),
    .sel (net2),
    .out (net348)
  );
  dff_cell flop112 (
    .d (net351),
    .clk (net1),
    .q (net350),
    .notq ()
  );
  mux_cell mux113 (
    .a (net352),
    .b (net353),
    .sel (net2),
    .out (net351)
  );
  dff_cell flop113 (
    .d (net354),
    .clk (net1),
    .q (net353),
    .notq ()
  );
  mux_cell mux114 (
    .a (net355),
    .b (net356),
    .sel (net2),
    .out (net354)
  );
  dff_cell flop114 (
    .d (net357),
    .clk (net1),
    .q (net356),
    .notq ()
  );
  mux_cell mux115 (
    .a (net358),
    .b (net359),
    .sel (net2),
    .out (net357)
  );
  dff_cell flop115 (
    .d (net360),
    .clk (net1),
    .q (net359),
    .notq ()
  );
  mux_cell mux116 (
    .a (net361),
    .b (net362),
    .sel (net2),
    .out (net360)
  );
  dff_cell flop116 (
    .d (net363),
    .clk (net1),
    .q (net362),
    .notq ()
  );
  mux_cell mux117 (
    .a (net364),
    .b (net365),
    .sel (net2),
    .out (net363)
  );
  dff_cell flop117 (
    .d (net366),
    .clk (net1),
    .q (net365),
    .notq ()
  );
  mux_cell mux118 (
    .a (net367),
    .b (net368),
    .sel (net2),
    .out (net366)
  );
  dff_cell flop118 (
    .d (net369),
    .clk (net1),
    .q (net368),
    .notq ()
  );
  mux_cell mux119 (
    .a (net370),
    .b (net371),
    .sel (net2),
    .out (net369)
  );
  dff_cell flop119 (
    .d (net372),
    .clk (net1),
    .q (net371),
    .notq ()
  );
  mux_cell mux120 (
    .a (net373),
    .b (net374),
    .sel (net2),
    .out (net372)
  );
  dff_cell flop120 (
    .d (net375),
    .clk (net1),
    .q (net374),
    .notq ()
  );
  mux_cell mux121 (
    .a (net376),
    .b (net377),
    .sel (net2),
    .out (net375)
  );
  dff_cell flop121 (
    .d (net378),
    .clk (net1),
    .q (net377),
    .notq ()
  );
  mux_cell mux122 (
    .a (net379),
    .b (net380),
    .sel (net2),
    .out (net378)
  );
  dff_cell flop122 (
    .d (net381),
    .clk (net1),
    .q (net380),
    .notq ()
  );
  mux_cell mux123 (
    .a (net382),
    .b (net383),
    .sel (net2),
    .out (net381)
  );
  dff_cell flop123 (
    .d (net385),
    .clk (net1),
    .q (net318),
    .notq ()
  );
  mux_cell mux124 (
    .a (net386),
    .b (net387),
    .sel (net2),
    .out (net385)
  );
  dff_cell flop124 (
    .d (net388),
    .clk (net1),
    .q (net387),
    .notq ()
  );
  mux_cell mux125 (
    .a (net389),
    .b (net390),
    .sel (net2),
    .out (net388)
  );
  dff_cell flop125 (
    .d (net391),
    .clk (net1),
    .q (net390),
    .notq ()
  );
  mux_cell mux126 (
    .a (net392),
    .b (net393),
    .sel (net2),
    .out (net391)
  );
  dff_cell flop126 (
    .d (net394),
    .clk (net1),
    .q (net393),
    .notq ()
  );
  mux_cell mux127 (
    .a (net395),
    .b (net333),
    .sel (net2),
    .out (net394)
  );
  dff_cell flop127 (
    .d (net396),
    .clk (net1),
    .q (net397),
    .notq ()
  );
  mux_cell mux128 (
    .a (net398),
    .b (net399),
    .sel (net2),
    .out (net396)
  );
  dff_cell flop128 (
    .d (net400),
    .clk (net1),
    .q (net399),
    .notq ()
  );
  mux_cell mux129 (
    .a (net401),
    .b (net402),
    .sel (net2),
    .out (net400)
  );
  dff_cell flop129 (
    .d (net403),
    .clk (net1),
    .q (net402),
    .notq ()
  );
  mux_cell mux130 (
    .a (net404),
    .b (net405),
    .sel (net2),
    .out (net403)
  );
  dff_cell flop130 (
    .d (net406),
    .clk (net1),
    .q (net405),
    .notq ()
  );
  mux_cell mux131 (
    .a (net407),
    .b (net408),
    .sel (net2),
    .out (net406)
  );
  dff_cell flop131 (
    .d (net409),
    .clk (net1),
    .q (net408),
    .notq ()
  );
  mux_cell mux132 (
    .a (net410),
    .b (net411),
    .sel (net2),
    .out (net409)
  );
  dff_cell flop132 (
    .d (net412),
    .clk (net1),
    .q (net411),
    .notq ()
  );
  mux_cell mux133 (
    .a (net413),
    .b (net414),
    .sel (net2),
    .out (net412)
  );
  dff_cell flop133 (
    .d (net415),
    .clk (net1),
    .q (net414),
    .notq ()
  );
  mux_cell mux134 (
    .a (net416),
    .b (net417),
    .sel (net2),
    .out (net415)
  );
  dff_cell flop134 (
    .d (net418),
    .clk (net1),
    .q (net417),
    .notq ()
  );
  mux_cell mux135 (
    .a (net419),
    .b (net420),
    .sel (net2),
    .out (net418)
  );
  dff_cell flop135 (
    .d (net421),
    .clk (net1),
    .q (net420),
    .notq ()
  );
  mux_cell mux136 (
    .a (net422),
    .b (net423),
    .sel (net2),
    .out (net421)
  );
  dff_cell flop136 (
    .d (net424),
    .clk (net1),
    .q (net423),
    .notq ()
  );
  mux_cell mux137 (
    .a (net425),
    .b (net426),
    .sel (net2),
    .out (net424)
  );
  dff_cell flop137 (
    .d (net427),
    .clk (net1),
    .q (net426),
    .notq ()
  );
  mux_cell mux138 (
    .a (net428),
    .b (net429),
    .sel (net2),
    .out (net427)
  );
  dff_cell flop138 (
    .d (net430),
    .clk (net1),
    .q (net429),
    .notq ()
  );
  mux_cell mux139 (
    .a (net431),
    .b (net432),
    .sel (net2),
    .out (net430)
  );
  dff_cell flop139 (
    .d (net433),
    .clk (net1),
    .q (net432),
    .notq ()
  );
  mux_cell mux140 (
    .a (net434),
    .b (net435),
    .sel (net2),
    .out (net433)
  );
  dff_cell flop140 (
    .d (net436),
    .clk (net1),
    .q (net435),
    .notq ()
  );
  mux_cell mux141 (
    .a (net437),
    .b (net438),
    .sel (net2),
    .out (net436)
  );
  dff_cell flop141 (
    .d (net439),
    .clk (net1),
    .q (net438),
    .notq ()
  );
  mux_cell mux142 (
    .a (net440),
    .b (net441),
    .sel (net2),
    .out (net439)
  );
  dff_cell flop142 (
    .d (net442),
    .clk (net1),
    .q (net441),
    .notq ()
  );
  mux_cell mux143 (
    .a (net443),
    .b (net444),
    .sel (net2),
    .out (net442)
  );
  dff_cell flop143 (
    .d (net445),
    .clk (net1),
    .q (net444),
    .notq ()
  );
  mux_cell mux144 (
    .a (net446),
    .b (net447),
    .sel (net2),
    .out (net445)
  );
  dff_cell flop144 (
    .d (net449),
    .clk (net1),
    .q (net383),
    .notq ()
  );
  mux_cell mux145 (
    .a (net450),
    .b (net451),
    .sel (net2),
    .out (net449)
  );
  dff_cell flop145 (
    .d (net452),
    .clk (net1),
    .q (net451),
    .notq ()
  );
  mux_cell mux146 (
    .a (net453),
    .b (net454),
    .sel (net2),
    .out (net452)
  );
  dff_cell flop146 (
    .d (net455),
    .clk (net1),
    .q (net454),
    .notq ()
  );
  mux_cell mux147 (
    .a (net456),
    .b (net457),
    .sel (net2),
    .out (net455)
  );
  dff_cell flop147 (
    .d (net458),
    .clk (net1),
    .q (net457),
    .notq ()
  );
  mux_cell mux148 (
    .a (net459),
    .b (net397),
    .sel (net2),
    .out (net458)
  );
  dff_cell flop148 (
    .d (net460),
    .clk (net1),
    .q (net461),
    .notq ()
  );
  mux_cell mux149 (
    .a (net462),
    .b (net463),
    .sel (net2),
    .out (net460)
  );
  dff_cell flop149 (
    .d (net464),
    .clk (net1),
    .q (net463),
    .notq ()
  );
  mux_cell mux150 (
    .a (net465),
    .b (net466),
    .sel (net2),
    .out (net464)
  );
  dff_cell flop150 (
    .d (net467),
    .clk (net1),
    .q (net466),
    .notq ()
  );
  mux_cell mux151 (
    .a (net468),
    .b (net469),
    .sel (net2),
    .out (net467)
  );
  dff_cell flop151 (
    .d (net470),
    .clk (net1),
    .q (net469),
    .notq ()
  );
  mux_cell mux152 (
    .a (net471),
    .b (net472),
    .sel (net2),
    .out (net470)
  );
  dff_cell flop152 (
    .d (net473),
    .clk (net1),
    .q (net472),
    .notq ()
  );
  mux_cell mux153 (
    .a (net474),
    .b (net475),
    .sel (net2),
    .out (net473)
  );
  dff_cell flop153 (
    .d (net476),
    .clk (net1),
    .q (net475),
    .notq ()
  );
  mux_cell mux154 (
    .a (net477),
    .b (net478),
    .sel (net2),
    .out (net476)
  );
  dff_cell flop154 (
    .d (net479),
    .clk (net1),
    .q (net478),
    .notq ()
  );
  mux_cell mux155 (
    .a (net480),
    .b (net481),
    .sel (net2),
    .out (net479)
  );
  dff_cell flop155 (
    .d (net482),
    .clk (net1),
    .q (net481),
    .notq ()
  );
  mux_cell mux156 (
    .a (net483),
    .b (net484),
    .sel (net2),
    .out (net482)
  );
  dff_cell flop156 (
    .d (net485),
    .clk (net1),
    .q (net484),
    .notq ()
  );
  mux_cell mux157 (
    .a (net486),
    .b (net487),
    .sel (net2),
    .out (net485)
  );
  dff_cell flop157 (
    .d (net488),
    .clk (net1),
    .q (net487),
    .notq ()
  );
  mux_cell mux158 (
    .a (net489),
    .b (net490),
    .sel (net2),
    .out (net488)
  );
  dff_cell flop158 (
    .d (net491),
    .clk (net1),
    .q (net490),
    .notq ()
  );
  mux_cell mux159 (
    .a (net492),
    .b (net493),
    .sel (net2),
    .out (net491)
  );
  dff_cell flop159 (
    .d (net494),
    .clk (net1),
    .q (net493),
    .notq ()
  );
  mux_cell mux160 (
    .a (net495),
    .b (net496),
    .sel (net2),
    .out (net494)
  );
  dff_cell flop160 (
    .d (net497),
    .clk (net1),
    .q (net496),
    .notq ()
  );
  mux_cell mux161 (
    .a (net498),
    .b (net499),
    .sel (net2),
    .out (net497)
  );
  dff_cell flop161 (
    .d (net500),
    .clk (net1),
    .q (net499),
    .notq ()
  );
  mux_cell mux162 (
    .a (net501),
    .b (net502),
    .sel (net2),
    .out (net500)
  );
  dff_cell flop162 (
    .d (net503),
    .clk (net1),
    .q (net502),
    .notq ()
  );
  mux_cell mux163 (
    .a (net504),
    .b (net505),
    .sel (net2),
    .out (net503)
  );
  dff_cell flop163 (
    .d (net506),
    .clk (net1),
    .q (net505),
    .notq ()
  );
  mux_cell mux164 (
    .a (net507),
    .b (net508),
    .sel (net2),
    .out (net506)
  );
  dff_cell flop164 (
    .d (net509),
    .clk (net1),
    .q (net508),
    .notq ()
  );
  mux_cell mux165 (
    .a (net510),
    .b (net4),
    .sel (net2),
    .out (net509)
  );
  dff_cell flop165 (
    .d (net512),
    .clk (net1),
    .q (net447),
    .notq ()
  );
  mux_cell mux166 (
    .a (net513),
    .b (net514),
    .sel (net2),
    .out (net512)
  );
  dff_cell flop166 (
    .d (net515),
    .clk (net1),
    .q (net514),
    .notq ()
  );
  mux_cell mux167 (
    .a (net516),
    .b (net517),
    .sel (net2),
    .out (net515)
  );
  dff_cell flop167 (
    .d (net518),
    .clk (net1),
    .q (net517),
    .notq ()
  );
  mux_cell mux168 (
    .a (net519),
    .b (net520),
    .sel (net2),
    .out (net518)
  );
  dff_cell flop168 (
    .d (net521),
    .clk (net1),
    .q (net520),
    .notq ()
  );
  mux_cell mux169 (
    .a (net522),
    .b (net461),
    .sel (net2),
    .out (net521)
  );
endmodule
