magic
tech sky130A
magscale 1 2
timestamp 1738411984
<< checkpaint >>
rect -1060 -1260 7832 7340
<< error_p >>
rect 6963 1833 6998 1867
rect 6964 1814 6998 1833
rect 6772 1765 6834 1771
rect 6772 1731 6784 1765
rect 6772 1725 6834 1731
rect 6772 437 6834 443
rect 6772 403 6784 437
rect 6772 397 6834 403
rect 6983 301 6998 1814
rect 7017 1780 7052 1814
rect 7372 1780 7407 1814
rect 7017 301 7051 1780
rect 7373 1761 7407 1780
rect 7181 1712 7243 1718
rect 7181 1678 7193 1712
rect 7181 1672 7243 1678
rect 7181 384 7243 390
rect 7181 350 7193 384
rect 7181 344 7243 350
rect 7017 267 7032 301
rect 7392 248 7407 1761
rect 7426 1727 7461 1761
rect 7426 248 7460 1727
rect 7590 1659 7652 1665
rect 7590 1625 7602 1659
rect 7590 1619 7652 1625
rect 7782 926 7816 944
rect 7782 890 7852 926
rect 7799 856 7870 890
rect 8150 856 8185 890
rect 7590 331 7652 337
rect 7590 297 7602 331
rect 7590 291 7652 297
rect 7426 214 7441 248
rect 7799 195 7869 856
rect 8151 837 8185 856
rect 7981 788 8039 794
rect 7981 754 7993 788
rect 7981 748 8039 754
rect 7981 278 8039 284
rect 7981 244 7993 278
rect 7981 238 8039 244
rect 7799 159 7852 195
rect 8170 142 8185 837
rect 8204 803 8239 837
rect 8519 803 8554 837
rect 8204 142 8238 803
rect 8520 784 8554 803
rect 8350 735 8408 741
rect 8350 701 8362 735
rect 8350 695 8408 701
rect 8350 225 8408 231
rect 8350 191 8362 225
rect 8350 185 8408 191
rect 8204 108 8219 142
rect 8539 89 8554 784
rect 8573 750 8608 784
rect 8573 89 8607 750
rect 8719 682 8777 688
rect 8719 648 8731 682
rect 8719 642 8777 648
rect 8719 172 8777 178
rect 8719 138 8731 172
rect 8719 132 8777 138
rect 8573 55 8588 89
use sky130_fd_pr__res_generic_l1_QHFG3U  R1
timestamp 1738407706
transform 1 0 100 0 1 300057
box -100 -300057 100 300057
use schmitt_trigger_ro  x1
timestamp 1738407706
transform 1 0 6625 0 1 318
box -53 -318 2334 1585
use sky130_fd_pr__cap_mim_m3_1_AHUHXA  XC1
timestamp 1738407706
transform 1 0 3386 0 1 3040
box -3186 -3040 3186 3040
<< end >>
