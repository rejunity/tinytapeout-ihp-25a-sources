magic
tech sky130A
magscale 1 2
timestamp 1741615844
<< nwell >>
rect 24423 3978 24784 4738
rect 25839 4636 28127 5183
rect 24539 3976 24722 3978
<< nmos >>
rect 24910 4560 24950 4660
rect 24910 4346 24950 4446
rect 25933 4353 25963 4553
rect 26020 4353 26050 4553
rect 24910 4052 24950 4252
rect 25010 4052 25210 4252
rect 25933 4099 25963 4299
rect 26220 4026 26300 4476
rect 26488 4353 26518 4553
rect 26575 4353 26605 4553
rect 26488 4099 26518 4299
rect 26775 4026 26855 4476
rect 27043 4353 27073 4553
rect 27130 4353 27160 4553
rect 27043 4099 27073 4299
rect 27330 4026 27410 4476
rect 27598 4353 27628 4553
rect 27685 4353 27715 4553
rect 27598 4099 27628 4299
rect 27885 4026 27965 4476
<< pmos >>
rect 25933 4926 25963 5126
rect 25933 4672 25963 4872
rect 26020 4672 26050 4872
rect 26220 4866 26290 5066
rect 26488 4926 26518 5126
rect 26488 4672 26518 4872
rect 26575 4672 26605 4872
rect 26775 4866 26845 5066
rect 27043 4926 27073 5126
rect 27043 4672 27073 4872
rect 27130 4672 27160 4872
rect 27330 4866 27400 5066
rect 27598 4926 27628 5126
rect 27598 4672 27628 4872
rect 27685 4672 27715 4872
rect 27885 4866 27955 5066
rect 24620 4496 24690 4596
rect 24620 4342 24690 4442
rect 24620 4014 24690 4214
<< ndiff >>
rect 24852 4648 24910 4660
rect 24852 4572 24864 4648
rect 24898 4572 24910 4648
rect 24852 4560 24910 4572
rect 24950 4648 25008 4660
rect 24950 4572 24962 4648
rect 24996 4572 25008 4648
rect 24950 4560 25008 4572
rect 24852 4434 24910 4446
rect 24852 4358 24864 4434
rect 24898 4358 24910 4434
rect 24852 4346 24910 4358
rect 24950 4434 25008 4446
rect 24950 4358 24962 4434
rect 24996 4358 25008 4434
rect 24950 4346 25008 4358
rect 24965 4252 24995 4346
rect 25875 4541 25933 4553
rect 25875 4365 25887 4541
rect 25921 4365 25933 4541
rect 25875 4353 25933 4365
rect 25963 4541 26020 4553
rect 25963 4365 25975 4541
rect 26009 4365 26020 4541
rect 25963 4353 26020 4365
rect 26050 4541 26108 4553
rect 26050 4365 26062 4541
rect 26096 4365 26108 4541
rect 26430 4541 26488 4553
rect 26050 4353 26108 4365
rect 26162 4464 26220 4476
rect 25875 4287 25933 4299
rect 24852 4240 24910 4252
rect 24852 4064 24864 4240
rect 24898 4064 24910 4240
rect 24852 4052 24910 4064
rect 24950 4052 25010 4252
rect 25210 4240 25268 4252
rect 25210 4064 25222 4240
rect 25256 4064 25268 4240
rect 25875 4111 25887 4287
rect 25921 4111 25933 4287
rect 25875 4099 25933 4111
rect 25963 4287 26021 4299
rect 25963 4111 25975 4287
rect 26009 4111 26021 4287
rect 25963 4099 26021 4111
rect 25210 4052 25268 4064
rect 26162 4038 26174 4464
rect 26208 4038 26220 4464
rect 26162 4026 26220 4038
rect 26300 4464 26358 4476
rect 26300 4038 26312 4464
rect 26346 4038 26358 4464
rect 26430 4365 26442 4541
rect 26476 4365 26488 4541
rect 26430 4353 26488 4365
rect 26518 4541 26575 4553
rect 26518 4365 26530 4541
rect 26564 4365 26575 4541
rect 26518 4353 26575 4365
rect 26605 4541 26663 4553
rect 26605 4365 26617 4541
rect 26651 4365 26663 4541
rect 26985 4541 27043 4553
rect 26605 4353 26663 4365
rect 26717 4464 26775 4476
rect 26430 4287 26488 4299
rect 26430 4111 26442 4287
rect 26476 4111 26488 4287
rect 26430 4099 26488 4111
rect 26518 4287 26576 4299
rect 26518 4111 26530 4287
rect 26564 4111 26576 4287
rect 26518 4099 26576 4111
rect 26300 4026 26358 4038
rect 26717 4038 26729 4464
rect 26763 4038 26775 4464
rect 26717 4026 26775 4038
rect 26855 4464 26913 4476
rect 26855 4038 26867 4464
rect 26901 4038 26913 4464
rect 26985 4365 26997 4541
rect 27031 4365 27043 4541
rect 26985 4353 27043 4365
rect 27073 4541 27130 4553
rect 27073 4365 27085 4541
rect 27119 4365 27130 4541
rect 27073 4353 27130 4365
rect 27160 4541 27218 4553
rect 27160 4365 27172 4541
rect 27206 4365 27218 4541
rect 27540 4541 27598 4553
rect 27160 4353 27218 4365
rect 27272 4464 27330 4476
rect 26985 4287 27043 4299
rect 26985 4111 26997 4287
rect 27031 4111 27043 4287
rect 26985 4099 27043 4111
rect 27073 4287 27131 4299
rect 27073 4111 27085 4287
rect 27119 4111 27131 4287
rect 27073 4099 27131 4111
rect 26855 4026 26913 4038
rect 27272 4038 27284 4464
rect 27318 4038 27330 4464
rect 27272 4026 27330 4038
rect 27410 4464 27468 4476
rect 27410 4038 27422 4464
rect 27456 4038 27468 4464
rect 27540 4365 27552 4541
rect 27586 4365 27598 4541
rect 27540 4353 27598 4365
rect 27628 4541 27685 4553
rect 27628 4365 27640 4541
rect 27674 4365 27685 4541
rect 27628 4353 27685 4365
rect 27715 4541 27773 4553
rect 27715 4365 27727 4541
rect 27761 4365 27773 4541
rect 27715 4353 27773 4365
rect 27827 4464 27885 4476
rect 27540 4287 27598 4299
rect 27540 4111 27552 4287
rect 27586 4111 27598 4287
rect 27540 4099 27598 4111
rect 27628 4287 27686 4299
rect 27628 4111 27640 4287
rect 27674 4111 27686 4287
rect 27628 4099 27686 4111
rect 27410 4026 27468 4038
rect 27827 4038 27839 4464
rect 27873 4038 27885 4464
rect 27827 4026 27885 4038
rect 27965 4464 28023 4476
rect 27965 4038 27977 4464
rect 28011 4038 28023 4464
rect 27965 4026 28023 4038
<< pdiff >>
rect 25875 5114 25933 5126
rect 25875 4938 25887 5114
rect 25921 4938 25933 5114
rect 25875 4926 25933 4938
rect 25963 5114 26021 5126
rect 25963 4938 25975 5114
rect 26009 4938 26021 5114
rect 26430 5114 26488 5126
rect 25963 4926 26021 4938
rect 26162 5054 26220 5066
rect 26162 4878 26174 5054
rect 26208 4878 26220 5054
rect 25875 4860 25933 4872
rect 25875 4684 25887 4860
rect 25921 4684 25933 4860
rect 25875 4672 25933 4684
rect 25963 4860 26020 4872
rect 25963 4684 25975 4860
rect 26009 4684 26020 4860
rect 25963 4672 26020 4684
rect 26050 4860 26108 4872
rect 26162 4866 26220 4878
rect 26290 5054 26348 5066
rect 26290 4878 26302 5054
rect 26336 4878 26348 5054
rect 26430 4938 26442 5114
rect 26476 4938 26488 5114
rect 26430 4926 26488 4938
rect 26518 5114 26576 5126
rect 26518 4938 26530 5114
rect 26564 4938 26576 5114
rect 26985 5114 27043 5126
rect 26518 4926 26576 4938
rect 26717 5054 26775 5066
rect 26290 4866 26348 4878
rect 26717 4878 26729 5054
rect 26763 4878 26775 5054
rect 26050 4684 26062 4860
rect 26096 4684 26108 4860
rect 26430 4860 26488 4872
rect 26050 4672 26108 4684
rect 26430 4684 26442 4860
rect 26476 4684 26488 4860
rect 26430 4672 26488 4684
rect 26518 4860 26575 4872
rect 26518 4684 26530 4860
rect 26564 4684 26575 4860
rect 26518 4672 26575 4684
rect 26605 4860 26663 4872
rect 26717 4866 26775 4878
rect 26845 5054 26903 5066
rect 26845 4878 26857 5054
rect 26891 4878 26903 5054
rect 26985 4938 26997 5114
rect 27031 4938 27043 5114
rect 26985 4926 27043 4938
rect 27073 5114 27131 5126
rect 27073 4938 27085 5114
rect 27119 4938 27131 5114
rect 27540 5114 27598 5126
rect 27073 4926 27131 4938
rect 27272 5054 27330 5066
rect 26845 4866 26903 4878
rect 27272 4878 27284 5054
rect 27318 4878 27330 5054
rect 26605 4684 26617 4860
rect 26651 4684 26663 4860
rect 26985 4860 27043 4872
rect 26605 4672 26663 4684
rect 26985 4684 26997 4860
rect 27031 4684 27043 4860
rect 26985 4672 27043 4684
rect 27073 4860 27130 4872
rect 27073 4684 27085 4860
rect 27119 4684 27130 4860
rect 27073 4672 27130 4684
rect 27160 4860 27218 4872
rect 27272 4866 27330 4878
rect 27400 5054 27458 5066
rect 27400 4878 27412 5054
rect 27446 4878 27458 5054
rect 27540 4938 27552 5114
rect 27586 4938 27598 5114
rect 27540 4926 27598 4938
rect 27628 5114 27686 5126
rect 27628 4938 27640 5114
rect 27674 4938 27686 5114
rect 27628 4926 27686 4938
rect 27827 5054 27885 5066
rect 27400 4866 27458 4878
rect 27827 4878 27839 5054
rect 27873 4878 27885 5054
rect 27160 4684 27172 4860
rect 27206 4684 27218 4860
rect 27540 4860 27598 4872
rect 27160 4672 27218 4684
rect 27540 4684 27552 4860
rect 27586 4684 27598 4860
rect 27540 4672 27598 4684
rect 27628 4860 27685 4872
rect 27628 4684 27640 4860
rect 27674 4684 27685 4860
rect 27628 4672 27685 4684
rect 27715 4860 27773 4872
rect 27827 4866 27885 4878
rect 27955 5054 28013 5066
rect 27955 4878 27967 5054
rect 28001 4878 28013 5054
rect 27955 4866 28013 4878
rect 27715 4684 27727 4860
rect 27761 4684 27773 4860
rect 27715 4672 27773 4684
rect 24562 4584 24620 4596
rect 24562 4508 24574 4584
rect 24608 4508 24620 4584
rect 24562 4496 24620 4508
rect 24690 4584 24748 4596
rect 24690 4508 24702 4584
rect 24736 4508 24748 4584
rect 24690 4496 24748 4508
rect 24562 4430 24620 4442
rect 24562 4354 24574 4430
rect 24608 4354 24620 4430
rect 24562 4342 24620 4354
rect 24690 4430 24748 4442
rect 24690 4354 24702 4430
rect 24736 4354 24748 4430
rect 24690 4342 24748 4354
rect 24562 4202 24620 4214
rect 24562 4026 24574 4202
rect 24608 4026 24620 4202
rect 24562 4014 24620 4026
rect 24690 4202 24748 4214
rect 24690 4026 24702 4202
rect 24736 4026 24748 4202
rect 24690 4014 24748 4026
<< ndiffc >>
rect 24864 4572 24898 4648
rect 24962 4572 24996 4648
rect 24864 4358 24898 4434
rect 24962 4358 24996 4434
rect 25887 4365 25921 4541
rect 25975 4365 26009 4541
rect 26062 4365 26096 4541
rect 24864 4064 24898 4240
rect 25222 4064 25256 4240
rect 25887 4111 25921 4287
rect 25975 4111 26009 4287
rect 26174 4038 26208 4464
rect 26312 4038 26346 4464
rect 26442 4365 26476 4541
rect 26530 4365 26564 4541
rect 26617 4365 26651 4541
rect 26442 4111 26476 4287
rect 26530 4111 26564 4287
rect 26729 4038 26763 4464
rect 26867 4038 26901 4464
rect 26997 4365 27031 4541
rect 27085 4365 27119 4541
rect 27172 4365 27206 4541
rect 26997 4111 27031 4287
rect 27085 4111 27119 4287
rect 27284 4038 27318 4464
rect 27422 4038 27456 4464
rect 27552 4365 27586 4541
rect 27640 4365 27674 4541
rect 27727 4365 27761 4541
rect 27552 4111 27586 4287
rect 27640 4111 27674 4287
rect 27839 4038 27873 4464
rect 27977 4038 28011 4464
<< pdiffc >>
rect 25887 4938 25921 5114
rect 25975 4938 26009 5114
rect 26174 4878 26208 5054
rect 25887 4684 25921 4860
rect 25975 4684 26009 4860
rect 26302 4878 26336 5054
rect 26442 4938 26476 5114
rect 26530 4938 26564 5114
rect 26729 4878 26763 5054
rect 26062 4684 26096 4860
rect 26442 4684 26476 4860
rect 26530 4684 26564 4860
rect 26857 4878 26891 5054
rect 26997 4938 27031 5114
rect 27085 4938 27119 5114
rect 27284 4878 27318 5054
rect 26617 4684 26651 4860
rect 26997 4684 27031 4860
rect 27085 4684 27119 4860
rect 27412 4878 27446 5054
rect 27552 4938 27586 5114
rect 27640 4938 27674 5114
rect 27839 4878 27873 5054
rect 27172 4684 27206 4860
rect 27552 4684 27586 4860
rect 27640 4684 27674 4860
rect 27967 4878 28001 5054
rect 27727 4684 27761 4860
rect 24574 4508 24608 4584
rect 24702 4508 24736 4584
rect 24574 4354 24608 4430
rect 24702 4354 24736 4430
rect 24574 4026 24608 4202
rect 24702 4026 24736 4202
<< psubdiff >>
rect 25212 4521 25262 4545
rect 25212 4345 25220 4521
rect 25254 4345 25262 4521
rect 25212 4321 25262 4345
rect 26202 3895 26348 3907
rect 26757 3895 26903 3907
rect 27312 3895 27458 3907
rect 27867 3895 28013 3907
rect 26191 3861 26215 3895
rect 26337 3861 26361 3895
rect 26746 3861 26770 3895
rect 26892 3861 26916 3895
rect 27301 3861 27325 3895
rect 27447 3861 27471 3895
rect 27856 3861 27880 3895
rect 28002 3861 28026 3895
rect 26202 3849 26348 3861
rect 26757 3849 26903 3861
rect 27312 3849 27458 3861
rect 27867 3849 28013 3861
<< nsubdiff >>
rect 26244 4796 26351 4808
rect 26233 4762 26257 4796
rect 26337 4762 26361 4796
rect 26244 4750 26351 4762
rect 26799 4796 26906 4808
rect 26788 4762 26812 4796
rect 26892 4762 26916 4796
rect 26799 4750 26906 4762
rect 27354 4796 27461 4808
rect 27343 4762 27367 4796
rect 27447 4762 27471 4796
rect 27354 4750 27461 4762
rect 27909 4796 28016 4808
rect 27898 4762 27922 4796
rect 28002 4762 28026 4796
rect 27909 4750 28016 4762
rect 24459 4304 24509 4328
rect 24459 4254 24467 4304
rect 24501 4254 24509 4304
rect 24459 4230 24509 4254
<< psubdiffcont >>
rect 25220 4345 25254 4521
rect 26215 3861 26337 3895
rect 26770 3861 26892 3895
rect 27325 3861 27447 3895
rect 27880 3861 28002 3895
<< nsubdiffcont >>
rect 26257 4762 26337 4796
rect 26812 4762 26892 4796
rect 27367 4762 27447 4796
rect 27922 4762 28002 4796
rect 24467 4254 24501 4304
<< poly >>
rect 25933 5126 25963 5152
rect 26220 5147 26290 5162
rect 26220 5113 26236 5147
rect 26274 5113 26290 5147
rect 26488 5126 26518 5152
rect 26775 5147 26845 5162
rect 26220 5066 26290 5113
rect 25933 4872 25963 4926
rect 26020 4872 26050 4898
rect 24620 4677 24690 4687
rect 24620 4643 24636 4677
rect 24674 4643 24690 4677
rect 24910 4660 24950 4686
rect 26775 5113 26791 5147
rect 26829 5113 26845 5147
rect 27043 5126 27073 5152
rect 27330 5147 27400 5162
rect 26775 5066 26845 5113
rect 26488 4872 26518 4926
rect 26575 4872 26605 4898
rect 26220 4840 26290 4866
rect 27330 5113 27346 5147
rect 27384 5113 27400 5147
rect 27598 5126 27628 5152
rect 27885 5147 27955 5162
rect 27330 5066 27400 5113
rect 27043 4872 27073 4926
rect 27130 4872 27160 4898
rect 26775 4840 26845 4866
rect 27885 5113 27901 5147
rect 27939 5113 27955 5147
rect 27885 5066 27955 5113
rect 27598 4872 27628 4926
rect 27685 4872 27715 4898
rect 27330 4840 27400 4866
rect 27885 4840 27955 4866
rect 24620 4596 24690 4643
rect 25759 4625 25825 4635
rect 25933 4625 25963 4672
rect 26020 4642 26050 4672
rect 25759 4591 25775 4625
rect 25809 4591 25963 4625
rect 25759 4581 25825 4591
rect 24910 4538 24950 4560
rect 25933 4553 25963 4591
rect 26005 4625 26070 4642
rect 26283 4625 26348 4641
rect 26488 4625 26518 4672
rect 26575 4642 26605 4672
rect 26005 4591 26020 4625
rect 26054 4591 26298 4625
rect 26332 4591 26518 4625
rect 26005 4575 26070 4591
rect 26283 4575 26348 4591
rect 26020 4553 26050 4575
rect 26488 4553 26518 4591
rect 26560 4625 26625 4642
rect 26838 4625 26903 4641
rect 27043 4625 27073 4672
rect 27130 4642 27160 4672
rect 26560 4591 26575 4625
rect 26609 4591 26853 4625
rect 26887 4591 27073 4625
rect 26560 4575 26625 4591
rect 26838 4575 26903 4591
rect 26575 4553 26605 4575
rect 27043 4553 27073 4591
rect 27115 4625 27180 4642
rect 27393 4625 27458 4641
rect 27598 4625 27628 4672
rect 27685 4642 27715 4672
rect 27115 4591 27130 4625
rect 27164 4591 27408 4625
rect 27442 4591 27628 4625
rect 27115 4575 27180 4591
rect 27393 4575 27458 4591
rect 27130 4553 27160 4575
rect 27598 4553 27628 4591
rect 27670 4625 27735 4642
rect 27948 4625 28013 4641
rect 27670 4591 27685 4625
rect 27719 4591 27963 4625
rect 27997 4591 28013 4625
rect 27670 4575 27735 4591
rect 27948 4575 28013 4591
rect 27685 4553 27715 4575
rect 24897 4522 24963 4538
rect 24620 4442 24690 4496
rect 24897 4488 24913 4522
rect 24947 4488 24963 4522
rect 24897 4472 24963 4488
rect 24910 4446 24950 4472
rect 24620 4295 24690 4342
rect 24910 4320 24950 4346
rect 24620 4261 24636 4295
rect 24674 4261 24690 4295
rect 24620 4214 24690 4261
rect 24910 4252 24950 4278
rect 26220 4476 26300 4502
rect 25933 4299 25963 4353
rect 26020 4327 26050 4353
rect 25010 4252 25210 4278
rect 25933 4073 25963 4099
rect 24910 4026 24950 4052
rect 25010 4026 25210 4052
rect 26775 4476 26855 4502
rect 26488 4299 26518 4353
rect 26575 4327 26605 4353
rect 26488 4073 26518 4099
rect 27330 4476 27410 4502
rect 27043 4299 27073 4353
rect 27130 4327 27160 4353
rect 27043 4073 27073 4099
rect 27885 4476 27965 4502
rect 27598 4299 27628 4353
rect 27685 4327 27715 4353
rect 27598 4073 27628 4099
rect 24910 4014 25210 4026
rect 24620 3988 24690 4014
rect 24910 3980 25045 4014
rect 25175 3980 25210 4014
rect 26220 4000 26300 4026
rect 26775 4000 26855 4026
rect 27330 4000 27410 4026
rect 27885 4000 27965 4026
rect 24910 3964 25210 3980
rect 26211 3988 26300 4000
rect 26211 3954 26227 3988
rect 26275 3954 26300 3988
rect 26211 3938 26300 3954
rect 26766 3988 26855 4000
rect 26766 3954 26782 3988
rect 26830 3954 26855 3988
rect 26766 3938 26855 3954
rect 27321 3988 27410 4000
rect 27321 3954 27337 3988
rect 27385 3954 27410 3988
rect 27321 3938 27410 3954
rect 27876 3988 27965 4000
rect 27876 3954 27892 3988
rect 27940 3954 27965 3988
rect 27876 3938 27965 3954
<< polycont >>
rect 26236 5113 26274 5147
rect 24636 4643 24674 4677
rect 26791 5113 26829 5147
rect 27346 5113 27384 5147
rect 27901 5113 27939 5147
rect 25775 4591 25809 4625
rect 26020 4591 26054 4625
rect 26298 4591 26332 4625
rect 26575 4591 26609 4625
rect 26853 4591 26887 4625
rect 27130 4591 27164 4625
rect 27408 4591 27442 4625
rect 27685 4591 27719 4625
rect 27963 4591 27997 4625
rect 24913 4488 24947 4522
rect 24636 4261 24674 4295
rect 25045 3980 25175 4014
rect 26227 3954 26275 3988
rect 26782 3954 26830 3988
rect 27337 3954 27385 3988
rect 27892 3954 27940 3988
<< locali >>
rect 25887 5164 26077 5198
rect 25887 5114 25921 5164
rect 25887 4922 25921 4938
rect 25975 5114 26009 5130
rect 26043 5070 26077 5164
rect 26442 5164 26632 5198
rect 26220 5113 26236 5147
rect 26274 5113 26290 5147
rect 26442 5114 26476 5164
rect 26043 5054 26208 5070
rect 26043 5036 26174 5054
rect 25975 4922 26009 4938
rect 25887 4860 25921 4876
rect 24620 4643 24636 4677
rect 24674 4643 24690 4677
rect 24864 4648 24898 4664
rect 24574 4584 24608 4600
rect 24574 4492 24608 4508
rect 24702 4584 24736 4600
rect 24864 4556 24898 4572
rect 24962 4648 24996 4664
rect 25775 4625 25809 4641
rect 25775 4575 25809 4591
rect 25887 4625 25921 4684
rect 25975 4860 26009 4876
rect 25975 4668 26009 4684
rect 26062 4860 26096 4876
rect 26174 4862 26208 4878
rect 26302 5054 26336 5070
rect 26442 4922 26476 4938
rect 26530 5114 26564 5130
rect 26598 5070 26632 5164
rect 26997 5164 27187 5198
rect 26775 5113 26791 5147
rect 26829 5113 26845 5147
rect 26997 5114 27031 5164
rect 26598 5054 26763 5070
rect 26598 5036 26729 5054
rect 26530 4922 26564 4938
rect 26302 4862 26336 4878
rect 26442 4860 26476 4876
rect 26233 4762 26257 4796
rect 26337 4762 26361 4796
rect 26096 4684 26208 4702
rect 26062 4668 26208 4684
rect 25887 4591 26020 4625
rect 26054 4591 26070 4625
rect 24962 4556 24996 4572
rect 25887 4541 25921 4591
rect 24702 4492 24736 4508
rect 24897 4488 24913 4522
rect 24947 4488 24963 4522
rect 25220 4521 25254 4537
rect 24574 4430 24608 4446
rect 24574 4338 24608 4354
rect 24702 4430 24736 4446
rect 24702 4338 24736 4354
rect 24864 4434 24898 4450
rect 24864 4342 24898 4358
rect 24962 4434 24996 4450
rect 24962 4342 24996 4358
rect 25887 4349 25921 4365
rect 25975 4541 26009 4557
rect 25975 4349 26009 4365
rect 26062 4541 26096 4557
rect 26062 4349 26096 4365
rect 26174 4464 26208 4668
rect 26442 4625 26476 4684
rect 26530 4860 26564 4876
rect 26530 4668 26564 4684
rect 26617 4860 26651 4876
rect 26729 4862 26763 4878
rect 26857 5054 26891 5070
rect 26997 4922 27031 4938
rect 27085 5114 27119 5130
rect 27153 5070 27187 5164
rect 27552 5164 27742 5198
rect 27330 5113 27346 5147
rect 27384 5113 27400 5147
rect 27552 5114 27586 5164
rect 27153 5054 27318 5070
rect 27153 5036 27284 5054
rect 27085 4922 27119 4938
rect 26857 4862 26891 4878
rect 26997 4860 27031 4876
rect 26788 4762 26812 4796
rect 26892 4762 26916 4796
rect 26651 4684 26763 4702
rect 26617 4668 26763 4684
rect 26282 4591 26298 4625
rect 26332 4591 26348 4625
rect 26442 4591 26575 4625
rect 26609 4591 26625 4625
rect 26442 4541 26476 4591
rect 25220 4329 25254 4345
rect 24467 4304 24501 4320
rect 24620 4261 24636 4295
rect 24674 4261 24690 4295
rect 25887 4287 25921 4303
rect 24467 4238 24501 4254
rect 24864 4240 24898 4256
rect 24574 4202 24608 4218
rect 24574 4010 24608 4026
rect 24702 4202 24736 4218
rect 24864 4048 24898 4064
rect 25222 4240 25256 4256
rect 25222 4048 25256 4064
rect 25887 4056 25921 4111
rect 25975 4287 26009 4303
rect 25975 4095 26009 4111
rect 24702 4010 24736 4026
rect 25887 4038 26174 4056
rect 25887 4022 26208 4038
rect 26312 4464 26346 4480
rect 26442 4349 26476 4365
rect 26530 4541 26564 4557
rect 26530 4349 26564 4365
rect 26617 4541 26651 4557
rect 26617 4349 26651 4365
rect 26729 4464 26763 4668
rect 26997 4625 27031 4684
rect 27085 4860 27119 4876
rect 27085 4668 27119 4684
rect 27172 4860 27206 4876
rect 27284 4862 27318 4878
rect 27412 5054 27446 5070
rect 27552 4922 27586 4938
rect 27640 5114 27674 5130
rect 27708 5070 27742 5164
rect 27885 5113 27901 5147
rect 27939 5113 27955 5147
rect 27708 5054 27873 5070
rect 27708 5036 27839 5054
rect 27640 4922 27674 4938
rect 27412 4862 27446 4878
rect 27552 4860 27586 4876
rect 27343 4762 27367 4796
rect 27447 4762 27471 4796
rect 27206 4684 27318 4702
rect 27172 4668 27318 4684
rect 26837 4591 26853 4625
rect 26887 4591 26903 4625
rect 26997 4591 27130 4625
rect 27164 4591 27180 4625
rect 26997 4541 27031 4591
rect 26312 4022 26346 4038
rect 26442 4287 26476 4303
rect 26442 4056 26476 4111
rect 26530 4287 26564 4303
rect 26530 4095 26564 4111
rect 26442 4038 26729 4056
rect 26442 4022 26763 4038
rect 26867 4464 26901 4480
rect 26997 4349 27031 4365
rect 27085 4541 27119 4557
rect 27085 4349 27119 4365
rect 27172 4541 27206 4557
rect 27172 4349 27206 4365
rect 27284 4464 27318 4668
rect 27552 4625 27586 4684
rect 27640 4860 27674 4876
rect 27640 4668 27674 4684
rect 27727 4860 27761 4876
rect 27839 4862 27873 4878
rect 27967 5054 28001 5070
rect 27967 4862 28001 4878
rect 27898 4762 27922 4796
rect 28002 4762 28026 4796
rect 27761 4684 27873 4702
rect 27727 4668 27873 4684
rect 27392 4591 27408 4625
rect 27442 4591 27458 4625
rect 27552 4591 27685 4625
rect 27719 4591 27735 4625
rect 27552 4541 27586 4591
rect 26867 4022 26901 4038
rect 26997 4287 27031 4303
rect 26997 4056 27031 4111
rect 27085 4287 27119 4303
rect 27085 4095 27119 4111
rect 26997 4038 27284 4056
rect 26997 4022 27318 4038
rect 27422 4464 27456 4480
rect 27552 4349 27586 4365
rect 27640 4541 27674 4557
rect 27640 4349 27674 4365
rect 27727 4541 27761 4557
rect 27727 4349 27761 4365
rect 27839 4464 27873 4668
rect 27947 4591 27963 4625
rect 27997 4591 28013 4625
rect 27422 4022 27456 4038
rect 27552 4287 27586 4303
rect 27552 4056 27586 4111
rect 27640 4287 27674 4303
rect 27640 4095 27674 4111
rect 27552 4038 27839 4056
rect 27552 4022 27873 4038
rect 27977 4464 28011 4480
rect 27977 4022 28011 4038
rect 25029 3980 25045 4014
rect 25175 3980 25191 4014
rect 25887 3741 25921 4022
rect 26211 3954 26227 3988
rect 26275 3954 26782 3988
rect 26830 3954 27337 3988
rect 27385 3954 27892 3988
rect 27940 3954 27965 3988
rect 26191 3861 26215 3895
rect 26337 3861 26361 3895
rect 26746 3861 26770 3895
rect 26892 3861 26916 3895
rect 27301 3861 27325 3895
rect 27447 3861 27471 3895
rect 27856 3861 27880 3895
rect 28002 3861 28026 3895
<< viali >>
rect 25887 4938 25921 5114
rect 25975 4938 26009 5114
rect 26236 5113 26274 5147
rect 26174 4878 26208 5054
rect 25887 4684 25921 4860
rect 24636 4643 24674 4677
rect 24574 4508 24608 4584
rect 24702 4508 24736 4584
rect 24864 4572 24898 4648
rect 24962 4572 24996 4648
rect 25775 4591 25809 4625
rect 25975 4684 26009 4860
rect 26302 4878 26336 5054
rect 26442 4938 26476 5114
rect 26530 4938 26564 5114
rect 26791 5113 26829 5147
rect 26729 4878 26763 5054
rect 26062 4684 26096 4860
rect 26257 4762 26337 4796
rect 26020 4591 26054 4625
rect 24913 4488 24947 4522
rect 24574 4354 24608 4430
rect 24702 4354 24736 4430
rect 24864 4358 24898 4434
rect 24962 4358 24996 4434
rect 25220 4345 25254 4521
rect 25887 4365 25921 4541
rect 25975 4365 26009 4541
rect 26062 4365 26096 4541
rect 26442 4684 26476 4860
rect 26530 4684 26564 4860
rect 26857 4878 26891 5054
rect 26997 4938 27031 5114
rect 27085 4938 27119 5114
rect 27346 5113 27384 5147
rect 27284 4878 27318 5054
rect 26617 4684 26651 4860
rect 26812 4762 26892 4796
rect 26298 4591 26332 4625
rect 26575 4591 26609 4625
rect 24467 4254 24501 4304
rect 24636 4261 24674 4295
rect 24574 4026 24608 4202
rect 24702 4026 24736 4202
rect 24864 4064 24898 4240
rect 25222 4064 25256 4240
rect 25887 4111 25921 4287
rect 25975 4111 26009 4287
rect 26174 4038 26208 4464
rect 26312 4038 26346 4464
rect 26442 4365 26476 4541
rect 26530 4365 26564 4541
rect 26617 4365 26651 4541
rect 26997 4684 27031 4860
rect 27085 4684 27119 4860
rect 27412 4878 27446 5054
rect 27552 4938 27586 5114
rect 27640 4938 27674 5114
rect 27901 5113 27939 5147
rect 27839 4878 27873 5054
rect 27172 4684 27206 4860
rect 27367 4762 27447 4796
rect 26853 4591 26887 4625
rect 27130 4591 27164 4625
rect 26442 4111 26476 4287
rect 26530 4111 26564 4287
rect 26729 4038 26763 4464
rect 26867 4038 26901 4464
rect 26997 4365 27031 4541
rect 27085 4365 27119 4541
rect 27172 4365 27206 4541
rect 27552 4684 27586 4860
rect 27640 4684 27674 4860
rect 27967 4878 28001 5054
rect 27727 4684 27761 4860
rect 27922 4762 28002 4796
rect 27408 4591 27442 4625
rect 27685 4591 27719 4625
rect 26997 4111 27031 4287
rect 27085 4111 27119 4287
rect 27284 4038 27318 4464
rect 27422 4038 27456 4464
rect 27552 4365 27586 4541
rect 27640 4365 27674 4541
rect 27727 4365 27761 4541
rect 27963 4591 27997 4625
rect 27552 4111 27586 4287
rect 27640 4111 27674 4287
rect 27839 4038 27873 4464
rect 27977 4038 28011 4464
rect 25045 3980 25175 4014
rect 26227 3954 26275 3988
rect 26782 3954 26830 3988
rect 27337 3954 27385 3988
rect 27892 3954 27940 3988
rect 26215 3861 26337 3895
rect 26770 3861 26892 3895
rect 27325 3861 27447 3895
rect 27880 3861 28002 3895
rect 25887 3707 25921 3741
<< metal1 >>
rect 25757 5165 27951 5198
rect 25757 5164 26841 5165
rect 25757 4832 25785 5164
rect 26220 5159 26841 5164
rect 26220 5147 26286 5159
rect 25881 5114 25927 5126
rect 25881 4938 25887 5114
rect 25921 4938 25927 5114
rect 25881 4926 25927 4938
rect 25969 5114 26015 5126
rect 25969 4938 25975 5114
rect 26009 4938 26015 5114
rect 26220 5113 26236 5147
rect 26274 5113 26286 5147
rect 26775 5147 26841 5159
rect 26220 5107 26286 5113
rect 26436 5114 26482 5126
rect 24640 4804 25785 4832
rect 25881 4860 25927 4872
rect 24640 4687 24668 4804
rect 24620 4677 24690 4687
rect 24620 4643 24636 4677
rect 24674 4643 24690 4677
rect 24620 4637 24690 4643
rect 24858 4648 24904 4660
rect 24568 4584 24614 4596
rect 24568 4508 24574 4584
rect 24608 4508 24614 4584
rect 24568 4496 24614 4508
rect 24696 4595 24742 4596
rect 24858 4595 24864 4648
rect 24696 4584 24864 4595
rect 24696 4508 24702 4584
rect 24736 4572 24864 4584
rect 24898 4572 24904 4648
rect 24736 4560 24904 4572
rect 24956 4659 25256 4687
rect 25881 4684 25887 4860
rect 25921 4684 25927 4860
rect 25881 4672 25927 4684
rect 25969 4860 26015 4938
rect 26168 5054 26214 5066
rect 26168 4878 26174 5054
rect 26208 4878 26214 5054
rect 26296 5054 26342 5066
rect 26296 4997 26302 5054
rect 26275 4991 26302 4997
rect 26275 4933 26302 4939
rect 25969 4684 25975 4860
rect 26009 4684 26015 4860
rect 25969 4672 26015 4684
rect 26056 4860 26102 4872
rect 26168 4866 26214 4878
rect 26296 4878 26302 4933
rect 26336 4878 26342 5054
rect 26436 4938 26442 5114
rect 26476 4938 26482 5114
rect 26436 4926 26482 4938
rect 26524 5114 26570 5126
rect 26524 4938 26530 5114
rect 26564 4938 26570 5114
rect 26775 5113 26791 5147
rect 26829 5113 26841 5147
rect 27330 5147 27396 5165
rect 26775 5107 26841 5113
rect 26991 5114 27037 5126
rect 26296 4866 26342 4878
rect 26056 4684 26062 4860
rect 26096 4684 26102 4860
rect 26056 4672 26102 4684
rect 24956 4648 25002 4659
rect 24956 4572 24962 4648
rect 24996 4572 25002 4648
rect 24956 4560 25002 4572
rect 24736 4549 24898 4560
rect 24736 4508 24742 4549
rect 24696 4496 24742 4508
rect 24864 4528 24898 4549
rect 25024 4531 25088 4537
rect 25024 4528 25030 4531
rect 24864 4522 25030 4528
rect 24277 4460 24341 4466
rect 24277 4408 24283 4460
rect 24335 4448 24341 4460
rect 24574 4448 24608 4496
rect 24864 4488 24913 4522
rect 24947 4488 25030 4522
rect 24864 4482 25030 4488
rect 25024 4479 25030 4482
rect 25082 4519 25088 4531
rect 25220 4527 25256 4659
rect 25757 4639 25785 4641
rect 25757 4633 25824 4639
rect 25757 4581 25766 4633
rect 25818 4581 25824 4633
rect 26005 4631 26070 4632
rect 26005 4625 26076 4631
rect 26005 4591 26020 4625
rect 26054 4591 26076 4625
rect 26005 4585 26076 4591
rect 25757 4575 25824 4581
rect 26174 4553 26208 4866
rect 26305 4802 26333 4866
rect 26436 4860 26482 4872
rect 26251 4796 26349 4802
rect 26245 4762 26257 4796
rect 26337 4762 26349 4796
rect 26251 4756 26349 4762
rect 26436 4684 26442 4860
rect 26476 4684 26482 4860
rect 26436 4672 26482 4684
rect 26524 4860 26570 4938
rect 26723 5054 26769 5066
rect 26723 4878 26729 5054
rect 26763 4878 26769 5054
rect 26851 5054 26897 5066
rect 26851 4997 26857 5054
rect 26835 4991 26857 4997
rect 26835 4933 26857 4939
rect 26524 4684 26530 4860
rect 26564 4684 26570 4860
rect 26524 4672 26570 4684
rect 26611 4860 26657 4872
rect 26723 4866 26769 4878
rect 26851 4878 26857 4933
rect 26891 4878 26897 5054
rect 26991 4938 26997 5114
rect 27031 4938 27037 5114
rect 26991 4926 27037 4938
rect 27079 5114 27125 5126
rect 27079 4938 27085 5114
rect 27119 4938 27125 5114
rect 27330 5113 27346 5147
rect 27384 5113 27396 5147
rect 27885 5147 27951 5165
rect 27330 5107 27396 5113
rect 27546 5114 27592 5126
rect 26851 4866 26897 4878
rect 26611 4684 26617 4860
rect 26651 4684 26657 4860
rect 26611 4672 26657 4684
rect 26283 4625 26408 4632
rect 26283 4591 26298 4625
rect 26332 4591 26408 4625
rect 26283 4585 26408 4591
rect 26560 4631 26625 4632
rect 26560 4625 26631 4631
rect 26560 4591 26575 4625
rect 26609 4591 26631 4625
rect 26560 4585 26631 4591
rect 25881 4541 25927 4553
rect 25214 4521 25260 4527
rect 25082 4491 25116 4519
rect 25082 4479 25088 4491
rect 25024 4473 25088 4479
rect 24335 4442 24608 4448
rect 24335 4430 24614 4442
rect 24335 4420 24574 4430
rect 24335 4408 24341 4420
rect 24277 4402 24341 4408
rect 24568 4354 24574 4420
rect 24608 4354 24614 4430
rect 24568 4342 24614 4354
rect 24696 4430 24742 4442
rect 24696 4354 24702 4430
rect 24736 4408 24742 4430
rect 24858 4434 24904 4446
rect 24858 4408 24864 4434
rect 24736 4380 24864 4408
rect 24736 4354 24742 4380
rect 24696 4342 24742 4354
rect 24858 4358 24864 4380
rect 24898 4358 24904 4434
rect 24858 4346 24904 4358
rect 24956 4434 25002 4446
rect 24956 4358 24962 4434
rect 24996 4358 25002 4434
rect 24956 4346 25002 4358
rect 25214 4345 25220 4521
rect 25254 4345 25260 4521
rect 25881 4365 25887 4541
rect 25921 4365 25927 4541
rect 25881 4353 25927 4365
rect 25969 4541 26015 4553
rect 25969 4365 25975 4541
rect 26009 4365 26015 4541
rect 24467 4310 24501 4320
rect 24461 4304 24507 4310
rect 24461 4254 24467 4304
rect 24501 4294 24507 4304
rect 24568 4294 24596 4342
rect 24702 4301 24736 4342
rect 25214 4339 25260 4345
rect 25220 4308 25256 4339
rect 24501 4266 24596 4294
rect 24501 4254 24507 4266
rect 24461 4248 24507 4254
rect 24465 4234 24501 4248
rect 24568 4214 24596 4266
rect 24624 4295 24736 4301
rect 24624 4261 24636 4295
rect 24674 4261 24736 4295
rect 24624 4255 24736 4261
rect 25168 4302 25256 4308
rect 24858 4240 24904 4252
rect 25220 4252 25256 4302
rect 25881 4287 25927 4299
rect 25220 4250 25262 4252
rect 25168 4244 25262 4250
rect 24568 4202 24614 4214
rect 24568 4026 24574 4202
rect 24608 4026 24614 4202
rect 24568 4014 24614 4026
rect 24696 4202 24742 4214
rect 24696 4026 24702 4202
rect 24736 4157 24742 4202
rect 24858 4157 24864 4240
rect 24736 4129 24864 4157
rect 24736 4026 24742 4129
rect 24696 4014 24742 4026
rect 24858 4064 24864 4129
rect 24898 4064 24904 4240
rect 24858 4020 24904 4064
rect 25215 4240 25262 4244
rect 25215 4064 25222 4240
rect 25256 4064 25262 4240
rect 25881 4111 25887 4287
rect 25921 4111 25927 4287
rect 25881 4099 25927 4111
rect 25969 4287 26015 4365
rect 26056 4541 26208 4553
rect 26056 4365 26062 4541
rect 26096 4515 26208 4541
rect 26096 4365 26102 4515
rect 26056 4353 26102 4365
rect 26168 4464 26214 4476
rect 25969 4111 25975 4287
rect 26009 4111 26015 4287
rect 25969 4099 26015 4111
rect 25215 4052 25262 4064
rect 26168 4038 26174 4464
rect 26208 4038 26214 4464
rect 26306 4464 26352 4476
rect 26306 4300 26312 4464
rect 26262 4248 26268 4300
rect 26168 4026 26214 4038
rect 26306 4038 26312 4248
rect 26346 4038 26352 4464
rect 26306 4026 26352 4038
rect 24858 4014 25187 4020
rect 24858 3980 25045 4014
rect 25175 3980 25187 4014
rect 25767 3997 25819 4003
rect 24858 3974 25187 3980
rect 25757 3953 25767 3989
rect 25819 3988 25857 3989
rect 26182 3988 26287 3994
rect 25819 3954 26227 3988
rect 26275 3954 26287 3988
rect 25819 3953 26287 3954
rect 26182 3948 26287 3953
rect 25767 3939 25819 3945
rect 26315 3901 26343 4026
rect 26380 4003 26408 4585
rect 26729 4553 26763 4866
rect 26860 4802 26888 4866
rect 26991 4860 27037 4872
rect 26806 4796 26904 4802
rect 26800 4762 26812 4796
rect 26892 4762 26904 4796
rect 26806 4756 26904 4762
rect 26991 4684 26997 4860
rect 27031 4684 27037 4860
rect 26991 4672 27037 4684
rect 27079 4860 27125 4938
rect 27278 5054 27324 5066
rect 27278 4878 27284 5054
rect 27318 4878 27324 5054
rect 27406 5054 27452 5066
rect 27406 4997 27412 5054
rect 27392 4991 27412 4997
rect 27392 4933 27412 4939
rect 27079 4684 27085 4860
rect 27119 4684 27125 4860
rect 27079 4672 27125 4684
rect 27166 4860 27212 4872
rect 27278 4866 27324 4878
rect 27406 4878 27412 4933
rect 27446 4878 27452 5054
rect 27546 4938 27552 5114
rect 27586 4938 27592 5114
rect 27546 4926 27592 4938
rect 27634 5114 27680 5126
rect 27634 4938 27640 5114
rect 27674 4938 27680 5114
rect 27885 5113 27901 5147
rect 27939 5113 27951 5147
rect 27885 5107 27951 5113
rect 27406 4866 27452 4878
rect 27166 4684 27172 4860
rect 27206 4684 27212 4860
rect 27166 4672 27212 4684
rect 26838 4625 26963 4632
rect 26838 4591 26853 4625
rect 26887 4591 26963 4625
rect 26838 4585 26963 4591
rect 27115 4631 27180 4632
rect 27115 4625 27186 4631
rect 27115 4591 27130 4625
rect 27164 4591 27186 4625
rect 27115 4585 27186 4591
rect 26436 4541 26482 4553
rect 26436 4365 26442 4541
rect 26476 4365 26482 4541
rect 26436 4353 26482 4365
rect 26524 4541 26570 4553
rect 26524 4365 26530 4541
rect 26564 4365 26570 4541
rect 26436 4287 26482 4299
rect 26436 4111 26442 4287
rect 26476 4111 26482 4287
rect 26436 4099 26482 4111
rect 26524 4287 26570 4365
rect 26611 4541 26763 4553
rect 26611 4365 26617 4541
rect 26651 4515 26763 4541
rect 26651 4365 26657 4515
rect 26611 4353 26657 4365
rect 26723 4464 26769 4476
rect 26524 4111 26530 4287
rect 26564 4111 26570 4287
rect 26524 4099 26570 4111
rect 26723 4038 26729 4464
rect 26763 4038 26769 4464
rect 26861 4464 26907 4476
rect 26861 4306 26867 4464
rect 26817 4300 26867 4306
rect 26817 4242 26867 4248
rect 26723 4026 26769 4038
rect 26861 4038 26867 4242
rect 26901 4038 26907 4464
rect 26861 4026 26907 4038
rect 26371 3997 26423 4003
rect 26737 3988 26842 3994
rect 26737 3954 26782 3988
rect 26830 3954 26842 3988
rect 26737 3948 26842 3954
rect 26371 3939 26423 3945
rect 26380 3938 26408 3939
rect 26870 3901 26898 4026
rect 26935 4003 26963 4585
rect 27284 4553 27318 4866
rect 27415 4802 27443 4866
rect 27546 4860 27592 4872
rect 27361 4796 27459 4802
rect 27355 4762 27367 4796
rect 27447 4762 27459 4796
rect 27361 4756 27459 4762
rect 27546 4684 27552 4860
rect 27586 4684 27592 4860
rect 27546 4672 27592 4684
rect 27634 4860 27680 4938
rect 27833 5054 27879 5066
rect 27833 4878 27839 5054
rect 27873 4878 27879 5054
rect 27961 5054 28007 5066
rect 27961 4991 27967 5054
rect 27932 4939 27938 4991
rect 27634 4684 27640 4860
rect 27674 4684 27680 4860
rect 27634 4672 27680 4684
rect 27721 4860 27767 4872
rect 27833 4866 27879 4878
rect 27961 4878 27967 4939
rect 28001 4878 28007 5054
rect 27961 4866 28007 4878
rect 27721 4684 27727 4860
rect 27761 4684 27767 4860
rect 27721 4672 27767 4684
rect 27393 4634 27457 4640
rect 27393 4582 27399 4634
rect 27451 4632 27457 4634
rect 27451 4585 27518 4632
rect 27670 4631 27735 4632
rect 27670 4625 27741 4631
rect 27670 4591 27685 4625
rect 27719 4591 27741 4625
rect 27670 4585 27741 4591
rect 27451 4582 27457 4585
rect 27393 4576 27457 4582
rect 26991 4541 27037 4553
rect 26991 4365 26997 4541
rect 27031 4365 27037 4541
rect 26991 4353 27037 4365
rect 27079 4541 27125 4553
rect 27079 4365 27085 4541
rect 27119 4365 27125 4541
rect 26991 4287 27037 4299
rect 26991 4111 26997 4287
rect 27031 4111 27037 4287
rect 26991 4099 27037 4111
rect 27079 4287 27125 4365
rect 27166 4541 27318 4553
rect 27166 4365 27172 4541
rect 27206 4515 27318 4541
rect 27206 4365 27212 4515
rect 27166 4353 27212 4365
rect 27278 4464 27324 4476
rect 27079 4111 27085 4287
rect 27119 4111 27125 4287
rect 27079 4099 27125 4111
rect 27278 4038 27284 4464
rect 27318 4038 27324 4464
rect 27416 4464 27462 4476
rect 27416 4306 27422 4464
rect 27392 4300 27422 4306
rect 27392 4242 27422 4248
rect 27278 4026 27324 4038
rect 27416 4038 27422 4242
rect 27456 4038 27462 4464
rect 27416 4026 27462 4038
rect 26926 3997 26978 4003
rect 27292 3988 27397 3994
rect 27292 3954 27337 3988
rect 27385 3954 27397 3988
rect 27292 3948 27397 3954
rect 26926 3939 26978 3945
rect 26935 3938 26966 3939
rect 27425 3901 27453 4026
rect 27490 4003 27518 4585
rect 27839 4553 27873 4866
rect 27970 4802 27998 4866
rect 27916 4796 28014 4802
rect 27910 4762 27922 4796
rect 28002 4762 28014 4796
rect 27916 4756 28014 4762
rect 27984 4632 28567 4633
rect 27948 4625 28567 4632
rect 27948 4591 27963 4625
rect 27997 4591 28567 4625
rect 27948 4585 28567 4591
rect 27546 4541 27592 4553
rect 27546 4365 27552 4541
rect 27586 4365 27592 4541
rect 27546 4353 27592 4365
rect 27634 4541 27680 4553
rect 27634 4365 27640 4541
rect 27674 4365 27680 4541
rect 27546 4287 27592 4299
rect 27546 4111 27552 4287
rect 27586 4111 27592 4287
rect 27546 4099 27592 4111
rect 27634 4287 27680 4365
rect 27721 4541 27873 4553
rect 27721 4365 27727 4541
rect 27761 4515 27873 4541
rect 27761 4365 27767 4515
rect 27721 4353 27767 4365
rect 27833 4464 27879 4476
rect 27634 4111 27640 4287
rect 27674 4111 27680 4287
rect 27634 4099 27680 4111
rect 27833 4038 27839 4464
rect 27873 4038 27879 4464
rect 27971 4464 28017 4476
rect 27971 4306 27977 4464
rect 27948 4300 27977 4306
rect 27948 4242 27977 4248
rect 27833 4026 27879 4038
rect 27971 4038 27977 4242
rect 28011 4038 28017 4464
rect 27971 4026 28017 4038
rect 27481 3997 27533 4003
rect 27847 3988 27952 3994
rect 27847 3954 27892 3988
rect 27940 3954 27952 3988
rect 27847 3948 27952 3954
rect 27481 3939 27533 3945
rect 27490 3938 27518 3939
rect 27980 3901 28008 4026
rect 26209 3895 26343 3901
rect 26764 3895 26898 3901
rect 27319 3895 27453 3901
rect 27874 3895 28008 3901
rect 26203 3861 26215 3895
rect 26337 3861 26349 3895
rect 26758 3861 26770 3895
rect 26892 3861 26904 3895
rect 27313 3861 27325 3895
rect 27447 3861 27459 3895
rect 27868 3861 27880 3895
rect 28002 3861 28014 3895
rect 26209 3855 26343 3861
rect 26764 3855 26898 3861
rect 27319 3855 27453 3861
rect 27874 3855 28008 3861
rect 28519 3796 28567 4585
rect 28519 3750 28568 3796
rect 25875 3741 25933 3747
rect 25875 3707 25887 3741
rect 25921 3707 25933 3741
rect 25875 3701 25933 3707
rect 25887 1483 25921 3701
rect 25887 1449 26621 1483
rect 26587 1038 26621 1449
rect 28520 1482 28568 3750
rect 28520 1434 30442 1482
rect 26498 894 26678 1038
rect 30394 984 30442 1434
rect 26492 714 26498 894
rect 26678 714 26684 894
rect 30362 732 30542 984
rect 30356 552 30362 732
rect 30542 552 30548 732
<< via1 >>
rect 26275 4939 26302 4991
rect 26302 4939 26327 4991
rect 24283 4408 24335 4460
rect 25030 4479 25082 4531
rect 25766 4625 25818 4633
rect 25766 4591 25775 4625
rect 25775 4591 25809 4625
rect 25809 4591 25818 4625
rect 25766 4581 25818 4591
rect 26835 4939 26857 4991
rect 26857 4939 26887 4991
rect 25168 4250 25220 4302
rect 26268 4248 26312 4300
rect 26312 4248 26320 4300
rect 25767 3945 25819 3997
rect 27392 4939 27412 4991
rect 27412 4939 27444 4991
rect 26817 4248 26867 4300
rect 26867 4248 26869 4300
rect 26371 3945 26423 3997
rect 27938 4939 27967 4991
rect 27967 4939 27990 4991
rect 27399 4625 27451 4634
rect 27399 4591 27408 4625
rect 27408 4591 27442 4625
rect 27442 4591 27451 4625
rect 27399 4582 27451 4591
rect 27392 4248 27422 4300
rect 27422 4248 27444 4300
rect 26926 3945 26978 3997
rect 27948 4248 27977 4300
rect 27977 4248 28000 4300
rect 27481 3945 27533 3997
rect 26498 714 26678 894
rect 30362 552 30542 732
<< metal2 >>
rect 27938 4991 27990 4997
rect 26269 4979 26275 4991
rect 24217 4951 26275 4979
rect 24217 4471 24245 4951
rect 26269 4939 26275 4951
rect 26327 4979 26333 4991
rect 26829 4979 26835 4991
rect 26327 4951 26835 4979
rect 26327 4939 26333 4951
rect 26829 4939 26835 4951
rect 26887 4979 26893 4991
rect 27386 4979 27392 4991
rect 26887 4951 27392 4979
rect 26887 4939 26893 4951
rect 27386 4939 27392 4951
rect 27444 4979 27450 4991
rect 27444 4951 27938 4979
rect 27444 4939 27450 4951
rect 27938 4933 27990 4939
rect 25760 4633 25824 4639
rect 25760 4581 25766 4633
rect 25818 4622 25824 4633
rect 27393 4634 27457 4640
rect 27393 4622 27399 4634
rect 25818 4594 27399 4622
rect 25818 4581 25824 4594
rect 25760 4575 25824 4581
rect 27393 4582 27399 4594
rect 27451 4582 27457 4634
rect 27393 4576 27457 4582
rect 25024 4531 25088 4537
rect 25024 4479 25030 4531
rect 25082 4519 25088 4531
rect 25082 4491 25296 4519
rect 25082 4479 25088 4491
rect 25024 4473 25088 4479
rect 24203 4466 24277 4471
rect 24203 4462 24341 4466
rect 24203 4406 24212 4462
rect 24268 4460 24341 4462
rect 24268 4408 24283 4460
rect 24335 4408 24341 4460
rect 24268 4406 24341 4408
rect 24203 4402 24341 4406
rect 24203 4397 24277 4402
rect 25053 4246 25062 4302
rect 25118 4288 25127 4302
rect 25162 4288 25168 4302
rect 25118 4260 25168 4288
rect 25118 4246 25127 4260
rect 25162 4250 25168 4260
rect 25220 4250 25226 4302
rect 25268 3985 25296 4491
rect 25324 4246 25333 4302
rect 25389 4288 25398 4302
rect 26268 4300 26320 4306
rect 25389 4260 26268 4288
rect 25389 4246 25398 4260
rect 26811 4288 26817 4300
rect 26320 4260 26817 4288
rect 26811 4248 26817 4260
rect 26869 4288 26875 4300
rect 27386 4288 27392 4300
rect 26869 4260 27392 4288
rect 26869 4248 26875 4260
rect 27386 4248 27392 4260
rect 27444 4288 27450 4300
rect 27942 4288 27948 4300
rect 27444 4260 27948 4288
rect 27444 4248 27450 4260
rect 27942 4248 27948 4260
rect 28000 4248 28006 4300
rect 26268 4242 26320 4248
rect 25761 3985 25767 3997
rect 25268 3957 25767 3985
rect 25761 3945 25767 3957
rect 25819 3945 25825 3997
rect 26365 3945 26371 3997
rect 26423 3945 26429 3997
rect 26920 3945 26926 3997
rect 26978 3945 26984 3997
rect 27475 3945 27481 3997
rect 27533 3988 27539 3997
rect 27533 3954 27762 3988
rect 27533 3945 27539 3954
rect 26383 3762 26411 3945
rect 26920 3939 26984 3945
rect 26938 3762 26966 3939
rect 27734 3762 27762 3954
rect 26360 3706 26369 3762
rect 26425 3706 26434 3762
rect 26915 3706 26924 3762
rect 26980 3706 26989 3762
rect 27711 3706 27720 3762
rect 27776 3706 27785 3762
rect 26498 894 26678 900
rect 26498 527 26678 714
rect 30362 732 30542 738
rect 26494 357 26503 527
rect 26673 357 26682 527
rect 30362 519 30542 552
rect 26498 352 26678 357
rect 30358 349 30367 519
rect 30537 349 30546 519
rect 30362 344 30542 349
<< via2 >>
rect 24212 4406 24268 4462
rect 25062 4246 25118 4302
rect 25333 4246 25389 4302
rect 26369 3706 26425 3762
rect 26924 3706 26980 3762
rect 27720 3706 27776 3762
rect 26503 357 26673 527
rect 30367 349 30537 519
<< metal3 >>
rect 410 4466 486 4472
rect 410 4402 416 4466
rect 480 4464 486 4466
rect 24203 4464 24273 4467
rect 480 4462 24273 4464
rect 480 4406 24212 4462
rect 24268 4406 24273 4462
rect 480 4404 24273 4406
rect 480 4402 486 4404
rect 410 4396 486 4402
rect 24203 4401 24273 4404
rect 24134 4242 24140 4306
rect 24204 4304 24210 4306
rect 25057 4304 25123 4307
rect 25328 4304 25394 4307
rect 24204 4302 25394 4304
rect 24204 4246 25062 4302
rect 25118 4246 25333 4302
rect 25389 4246 25394 4302
rect 24204 4244 25394 4246
rect 24204 4242 24210 4244
rect 25057 4241 25123 4244
rect 25328 4241 25394 4244
rect 25756 4076 26412 5264
rect 25756 4008 26427 4076
rect 26667 4018 27323 5274
rect 26367 3767 26427 4008
rect 26922 3767 26982 4018
rect 27563 4008 28219 5264
rect 27718 3767 27778 4008
rect 26364 3762 26430 3767
rect 26364 3706 26369 3762
rect 26425 3706 26430 3762
rect 26364 3701 26430 3706
rect 26919 3762 26985 3767
rect 26919 3706 26924 3762
rect 26980 3706 26985 3762
rect 26919 3701 26985 3706
rect 27715 3762 27781 3767
rect 27715 3706 27720 3762
rect 27776 3706 27781 3762
rect 27715 3701 27781 3706
rect 26498 527 26678 532
rect 26498 357 26503 527
rect 26673 357 26678 527
rect 26498 213 26678 357
rect 26498 172 26562 213
rect 26556 149 26562 172
rect 26626 172 26678 213
rect 30362 519 30542 524
rect 30362 349 30367 519
rect 30537 349 30542 519
rect 30362 220 30542 349
rect 30362 198 30410 220
rect 26626 149 26632 172
rect 30404 156 30410 198
rect 30474 198 30542 220
rect 30474 156 30480 198
rect 30404 150 30480 156
rect 26556 143 26632 149
<< via3 >>
rect 416 4402 480 4466
rect 24140 4242 24204 4306
rect 26562 149 26626 213
rect 30410 156 30474 220
<< mimcap >>
rect 25784 5196 26384 5236
rect 25784 4076 25824 5196
rect 26344 4076 26384 5196
rect 25784 4036 26384 4076
rect 26695 5206 27295 5246
rect 26695 4086 26735 5206
rect 27255 4086 27295 5206
rect 26695 4046 27295 4086
rect 27591 5196 28191 5236
rect 27591 4076 27631 5196
rect 28151 4076 28191 5196
rect 27591 4036 28191 4076
<< mimcapcontact >>
rect 25824 4076 26344 5196
rect 26735 4086 27255 5206
rect 27631 4076 28151 5196
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 4466 600 44152
rect 200 4402 416 4466
rect 480 4402 600 4466
rect 200 1000 600 4402
rect 800 4304 1200 44152
rect 26734 5206 27256 5207
rect 25823 5196 26345 5197
rect 25823 5057 25824 5196
rect 24139 4996 25824 5057
rect 24139 4307 24200 4996
rect 24139 4306 24205 4307
rect 24139 4304 24140 4306
rect 800 4244 24140 4304
rect 800 1000 1200 4244
rect 24139 4242 24140 4244
rect 24204 4242 24205 4306
rect 24139 4241 24205 4242
rect 25823 4076 25824 4996
rect 26344 5057 26345 5196
rect 26734 5057 26735 5206
rect 26344 4997 26735 5057
rect 26344 4076 26345 4997
rect 26734 4086 26735 4997
rect 27255 5057 27256 5206
rect 27630 5196 28152 5197
rect 27630 5057 27631 5196
rect 27255 4997 27631 5057
rect 27255 4086 27256 4997
rect 26734 4085 27256 4086
rect 25823 4075 26345 4076
rect 27630 4076 27631 4997
rect 28151 4076 28152 5196
rect 27630 4075 28152 4076
rect 30404 220 30480 226
rect 26556 213 26632 219
rect 26556 200 26562 213
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 149 26562 200
rect 26626 200 26632 213
rect 30404 200 30410 220
rect 26626 149 26678 200
rect 26498 0 26678 149
rect 30362 156 30410 200
rect 30474 200 30480 220
rect 30474 156 30542 200
rect 30362 0 30542 156
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal2 25082 4491 25116 4519 3 bias.Vnbias
rlabel metal1 24620 4637 24690 4687 1 bias.Vpbias
rlabel metal1 25220 4240 25249 4687 3 bias.VSS
rlabel metal1 24568 4014 24614 4015 5 bias.VDD
<< end >>
