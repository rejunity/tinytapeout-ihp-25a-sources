/* Automatically generated from https://wokwi.com/projects/413387190167208961 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_413387190167208961(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = ui_in[0];
  wire net2 = ui_in[1];
  wire net3 = ui_in[2];
  wire net4 = ui_in[3];
  wire net5 = ui_in[4];
  wire net6 = ui_in[5];
  wire net7 = ui_in[6];
  wire net8 = ui_in[7];
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13 = 1'b0;
  wire net14 = 1'b0;
  wire net15 = 1'b1;
  wire net16 = 1'b1;
  wire net17 = 1'b0;
  wire net18 = 1'b1;

  assign uo_out[0] = net9;
  assign uo_out[1] = net10;
  assign uo_out[2] = net11;
  assign uo_out[3] = net12;
  assign uo_out[4] = 0;
  assign uo_out[5] = 0;
  assign uo_out[6] = 0;
  assign uo_out[7] = 0;
  assign uio_out[0] = net13;
  assign uio_oe[0] = net13;
  assign uio_out[1] = net13;
  assign uio_oe[1] = net13;
  assign uio_out[2] = net13;
  assign uio_oe[2] = net13;
  assign uio_out[3] = net13;
  assign uio_oe[3] = net13;
  assign uio_out[4] = net14;
  assign uio_oe[4] = net14;
  assign uio_out[5] = net14;
  assign uio_oe[5] = net14;
  assign uio_out[6] = net14;
  assign uio_oe[6] = net14;
  assign uio_out[7] = net14;
  assign uio_oe[7] = net14;

  nand_cell nand1 (
    .a (net7),
    .b (net8),
    .out (net12)
  );
  nand_cell nand5 (
    .a (net5),
    .b (net6),
    .out (net11)
  );
  nand_cell nand6 (
    .a (net3),
    .b (net4),
    .out (net10)
  );
  nand_cell nand7 (
    .a (net1),
    .b (net2),
    .out (net9)
  );
endmodule
