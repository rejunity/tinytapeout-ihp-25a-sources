** sch_path: /foss/designs/tt10-uR-IPs/xschem/T1/schmTrigg/schmTrigg.sch
.subckt schmTrigg Vin VSS VDD Vout
*.PININFO Vin:I VDD:I VSS:I Vout:O
XM1 VDD Vout Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Vn Vin VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 Vout Vin Vn Vn sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 VSS Vout Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 Vout Vin Vp Vp sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Vp Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
