magic
tech sky130A
magscale 1 2
timestamp 1738407706
<< error_s >>
rect 338 1515 373 1549
rect 339 1496 373 1515
rect 147 1447 209 1453
rect 147 1413 159 1447
rect 147 1407 209 1413
rect 147 119 209 125
rect 147 85 159 119
rect 147 79 209 85
rect 358 -17 373 1496
rect 392 1462 427 1496
rect 747 1462 782 1496
rect 392 -17 426 1462
rect 748 1443 782 1462
rect 556 1394 618 1400
rect 556 1360 568 1394
rect 556 1354 618 1360
rect 556 66 618 72
rect 556 32 568 66
rect 556 26 618 32
rect 392 -51 407 -17
rect 767 -70 782 1443
rect 801 1409 836 1443
rect 801 -70 835 1409
rect 965 1341 1027 1347
rect 965 1307 977 1341
rect 965 1301 1027 1307
rect 1157 608 1191 626
rect 1157 572 1227 608
rect 1174 538 1245 572
rect 1525 538 1560 572
rect 965 13 1027 19
rect 965 -21 977 13
rect 965 -27 1027 -21
rect 801 -104 816 -70
rect 1174 -123 1244 538
rect 1526 519 1560 538
rect 1356 470 1414 476
rect 1356 436 1368 470
rect 1356 430 1414 436
rect 1356 -40 1414 -34
rect 1356 -74 1368 -40
rect 1356 -80 1414 -74
rect 1174 -159 1227 -123
rect 1545 -176 1560 519
rect 1579 485 1614 519
rect 1894 485 1929 519
rect 1579 -176 1613 485
rect 1895 466 1929 485
rect 1725 417 1783 423
rect 1725 383 1737 417
rect 1725 377 1783 383
rect 1725 -93 1783 -87
rect 1725 -127 1737 -93
rect 1725 -133 1783 -127
rect 1579 -210 1594 -176
rect 1914 -229 1929 466
rect 1948 432 1983 466
rect 1948 -229 1982 432
rect 2094 364 2152 370
rect 2094 330 2106 364
rect 2094 324 2152 330
rect 2094 -146 2152 -140
rect 2094 -180 2106 -146
rect 2094 -186 2152 -180
rect 1948 -263 1963 -229
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM1
timestamp 1738407706
transform 1 0 1754 0 1 145
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM2
timestamp 1738407706
transform 1 0 587 0 1 713
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM3
timestamp 1738407706
transform 1 0 2123 0 1 92
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM4
timestamp 1738407706
transform 1 0 996 0 1 660
box -231 -819 231 819
use sky130_fd_pr__nfet_01v8_lvt_UH8C49  XM6
timestamp 1738407706
transform 1 0 1385 0 1 198
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_MT5C5V  XM10
timestamp 1738407706
transform 1 0 178 0 1 766
box -231 -819 231 819
<< end >>
