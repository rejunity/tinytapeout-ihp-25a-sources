magic
tech sky130A
magscale 1 2
timestamp 1741560270
<< error_p >>
rect -98 -194 -40 256
rect 40 -194 98 256
rect -45 -232 27 -226
rect -45 -266 -33 -232
rect -45 -272 27 -266
<< nmos >>
rect -40 -194 40 256
<< ndiff >>
rect -98 244 -40 256
rect -98 -182 -86 244
rect -52 -182 -40 244
rect -98 -194 -40 -182
rect 40 244 98 256
rect 40 -182 52 244
rect 86 -182 98 244
rect 40 -194 98 -182
<< ndiffc >>
rect -86 -182 -52 244
rect 52 -182 86 244
<< poly >>
rect -40 256 40 282
rect -40 -220 40 -194
rect -49 -232 40 -220
rect -49 -266 -33 -232
rect 15 -266 40 -232
rect -49 -282 40 -266
<< polycont >>
rect -33 -266 15 -232
<< locali >>
rect -86 244 -52 260
rect -86 -198 -52 -182
rect 52 244 86 260
rect 52 -198 86 -182
rect -49 -266 -33 -232
rect 15 -266 31 -232
<< viali >>
rect -86 -182 -52 244
rect 52 -182 86 244
rect -33 -266 15 -232
<< metal1 >>
rect -92 244 -46 256
rect -92 -182 -86 244
rect -52 -182 -46 244
rect -92 -194 -46 -182
rect 46 244 92 256
rect 46 -182 52 244
rect 86 -182 92 244
rect 46 -194 92 -182
rect -45 -232 27 -226
rect -45 -266 -33 -232
rect 15 -266 27 -232
rect -45 -272 27 -266
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.25 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
