magic
tech sky130A
magscale 1 2
timestamp 1741535882
<< metal3 >>
rect -474 -328 182 328
<< mimcap >>
rect -446 260 154 300
rect -446 -260 -406 260
rect 114 -260 154 260
rect -446 -300 154 -260
<< mimcapcontact >>
rect -406 -260 114 260
<< metal4 >>
rect -407 260 115 261
rect -407 -260 -406 260
rect 114 -260 115 260
rect -407 -261 115 -260
<< properties >>
string FIXED_BBOX -486 -340 194 340
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3 l 3 val 20.28 carea 2.00 cperi 0.19 class capacitor nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
