/* Automatically generated from https://wokwi.com/projects/414123795172381697 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_414123795172381697(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = rst_n;
  wire net3 = ui_in[0];
  wire net4 = ui_in[1];
  wire net5 = ui_in[2];
  wire net6 = ui_in[3];
  wire net7 = ui_in[4];
  wire net8 = ui_in[5];
  wire net9 = ui_in[6];
  wire net10 = ui_in[7];
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18 = 1'b0;
  wire net19 = 1'b1;
  wire net20 = 1'b1;
  wire net21 = 1'b0;
  wire net22 = 1'b1;
  wire net23;
  wire net24 = 1'b0;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35 = 1'b0;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49 = 1'b0;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103 = 1'b0;
  wire net104;
  wire net105;
  wire net106;
  wire net107 = 1'b1;
  wire net108;
  wire net109 = 1'b0;
  wire net110;
  wire net111;
  wire net112;
  wire net113 = 1'b0;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118 = 1'b0;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123 = 1'b0;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128 = 1'b0;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134 = 1'b0;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139 = 1'b0;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144 = 1'b0;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149 = 1'b0;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154 = 1'b0;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159 = 1'b0;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164 = 1'b0;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169 = 1'b0;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174 = 1'b0;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179 = 1'b0;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208 = 1'b0;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213 = 1'b0;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225 = 1'b0;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230 = 1'b0;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;

  assign uo_out[0] = net11;
  assign uo_out[1] = net12;
  assign uo_out[2] = net13;
  assign uo_out[3] = net14;
  assign uo_out[4] = net15;
  assign uo_out[5] = net16;
  assign uo_out[6] = net17;
  assign uo_out[7] = 0;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  dffsr_cell flop1 (
    .d (net23),
    .clk (net1),
    .s (net24),
    .r (net25),
    .q (net26),
    .notq (net27)
  );
  dffsr_cell flop2 (
    .d (net28),
    .clk (net1),
    .s (net24),
    .r (net25),
    .q (net29),
    .notq (net30)
  );
  dffsr_cell flop3 (
    .d (net31),
    .clk (net1),
    .s (net24),
    .r (net25),
    .q (net32),
    .notq (net33)
  );
  dffsr_cell flop4 (
    .d (net34),
    .clk (net1),
    .s (net25),
    .r (net35),
    .q (net36),
    .notq (net37)
  );
  dffsr_cell flop5 (
    .d (net38),
    .clk (net1),
    .s (net35),
    .r (net25),
    .q (net39),
    .notq (net40)
  );
  dffsr_cell flop6 (
    .d (net41),
    .clk (net1),
    .s (net25),
    .r (net35),
    .q (net42),
    .notq (net43)
  );
  mux_cell mux1 (
    .a (net23),
    .b (net44),
    .sel (net45),
    .out (net23)
  );
  mux_cell mux2 (
    .a (net28),
    .b (net46),
    .sel (net45),
    .out (net28)
  );
  mux_cell mux3 (
    .a (net31),
    .b (net47),
    .sel (net45),
    .out (net31)
  );
  mux_cell mux4 (
    .a (net34),
    .b (net26),
    .sel (net45),
    .out (net34)
  );
  mux_cell mux5 (
    .a (net38),
    .b (net29),
    .sel (net45),
    .out (net38)
  );
  mux_cell mux6 (
    .a (net41),
    .b (net32),
    .sel (net45),
    .out (net41)
  );
  dffsr_cell flop7 (
    .d (net48),
    .clk (net1),
    .s (net49),
    .r (net25),
    .q (net50),
    .notq (net51)
  );
  dffsr_cell flop8 (
    .d (net52),
    .clk (net1),
    .s (net49),
    .r (net25),
    .q (net53),
    .notq (net54)
  );
  dffsr_cell flop9 (
    .d (net55),
    .clk (net1),
    .s (net25),
    .r (net49),
    .q (net56),
    .notq (net57)
  );
  mux_cell mux7 (
    .a (net48),
    .b (net36),
    .sel (net45),
    .out (net48)
  );
  mux_cell mux8 (
    .a (net52),
    .b (net39),
    .sel (net45),
    .out (net52)
  );
  mux_cell mux9 (
    .a (net55),
    .b (net42),
    .sel (net45),
    .out (net55)
  );
  not_cell not5 (
    .in (net2),
    .out (net25)
  );
  and_cell and1 (
    .a (net33),
    .b (net30),
    .out (net58)
  );
  and_cell and2 (
    .a (net27),
    .b (net58),
    .out (net59)
  );
  and_cell and3 (
    .a (net26),
    .b (net58),
    .out (net60)
  );
  and_cell and4 (
    .a (net33),
    .b (net29),
    .out (net61)
  );
  and_cell and5 (
    .a (net27),
    .b (net61),
    .out (net62)
  );
  and_cell and6 (
    .a (net26),
    .b (net61),
    .out (net63)
  );
  and_cell and7 (
    .a (net27),
    .b (net64),
    .out (net65)
  );
  and_cell and8 (
    .a (net26),
    .b (net64),
    .out (net66)
  );
  and_cell and9 (
    .a (net29),
    .b (net32),
    .out (net67)
  );
  and_cell and10 (
    .a (net30),
    .b (net32),
    .out (net64)
  );
  and_cell and11 (
    .a (net43),
    .b (net40),
    .out (net68)
  );
  and_cell and12 (
    .a (net37),
    .b (net68),
    .out (net69)
  );
  and_cell and13 (
    .a (net36),
    .b (net68),
    .out (net70)
  );
  and_cell and14 (
    .a (net43),
    .b (net39),
    .out (net71)
  );
  and_cell and15 (
    .a (net37),
    .b (net71),
    .out (net72)
  );
  and_cell and16 (
    .a (net36),
    .b (net71),
    .out (net73)
  );
  and_cell and17 (
    .a (net37),
    .b (net74),
    .out (net75)
  );
  and_cell and18 (
    .a (net36),
    .b (net74),
    .out (net76)
  );
  and_cell and19 (
    .a (net39),
    .b (net42),
    .out (net77)
  );
  and_cell and20 (
    .a (net40),
    .b (net42),
    .out (net74)
  );
  and_cell and21 (
    .a (net57),
    .b (net54),
    .out (net78)
  );
  and_cell and22 (
    .a (net51),
    .b (net78),
    .out (net79)
  );
  and_cell and23 (
    .a (net50),
    .b (net78),
    .out (net80)
  );
  and_cell and24 (
    .a (net57),
    .b (net53),
    .out (net81)
  );
  and_cell and25 (
    .a (net51),
    .b (net81),
    .out (net82)
  );
  and_cell and26 (
    .a (net50),
    .b (net81),
    .out (net83)
  );
  and_cell and27 (
    .a (net51),
    .b (net84),
    .out (net85)
  );
  and_cell and28 (
    .a (net50),
    .b (net84),
    .out (net86)
  );
  and_cell and29 (
    .a (net53),
    .b (net56),
    .out (net87)
  );
  and_cell and30 (
    .a (net54),
    .b (net56),
    .out (net84)
  );
  or_cell or3 (
    .a (net69),
    .b (net79),
    .out (net88)
  );
  or_cell or4 (
    .a (net70),
    .b (net80),
    .out (net89)
  );
  or_cell or5 (
    .a (net72),
    .b (net82),
    .out (net90)
  );
  or_cell or6 (
    .a (net73),
    .b (net83),
    .out (net91)
  );
  or_cell or7 (
    .a (net75),
    .b (net85),
    .out (net92)
  );
  or_cell or8 (
    .a (net76),
    .b (net86),
    .out (net93)
  );
  or_cell or9 (
    .a (net77),
    .b (net87),
    .out (net94)
  );
  or_cell or2 (
    .a (net59),
    .b (net88),
    .out (net95)
  );
  or_cell or10 (
    .a (net60),
    .b (net89),
    .out (net96)
  );
  or_cell or11 (
    .a (net62),
    .b (net90),
    .out (net97)
  );
  or_cell or12 (
    .a (net63),
    .b (net91),
    .out (net98)
  );
  or_cell or13 (
    .a (net65),
    .b (net92),
    .out (net99)
  );
  or_cell or14 (
    .a (net66),
    .b (net93),
    .out (net100)
  );
  or_cell or15 (
    .a (net67),
    .b (net94),
    .out (net101)
  );
  dffsr_cell flop10 (
    .d (net102),
    .clk (net1),
    .s (net103),
    .r (net104),
    .q (net105),
    .notq (net106)
  );
  mux_cell mux10 (
    .a (net105),
    .b (net106),
    .sel (net107),
    .out (net102)
  );
  dffsr_cell flop11 (
    .d (net108),
    .clk (net1),
    .s (net109),
    .r (net104),
    .q (net110),
    .notq (net111)
  );
  mux_cell mux11 (
    .a (net110),
    .b (net111),
    .sel (net105),
    .out (net108)
  );
  dffsr_cell flop12 (
    .d (net112),
    .clk (net1),
    .s (net113),
    .r (net104),
    .q (net114),
    .notq (net115)
  );
  mux_cell mux12 (
    .a (net114),
    .b (net115),
    .sel (net116),
    .out (net112)
  );
  and_cell and31 (
    .a (net110),
    .b (net105),
    .out (net116)
  );
  dffsr_cell flop13 (
    .d (net117),
    .clk (net1),
    .s (net118),
    .r (net104),
    .q (net119),
    .notq (net120)
  );
  mux_cell mux13 (
    .a (net119),
    .b (net120),
    .sel (net121),
    .out (net117)
  );
  and_cell and32 (
    .a (net114),
    .b (net116),
    .out (net121)
  );
  dffsr_cell flop14 (
    .d (net122),
    .clk (net1),
    .s (net123),
    .r (net104),
    .q (net124),
    .notq (net125)
  );
  mux_cell mux14 (
    .a (net124),
    .b (net125),
    .sel (net126),
    .out (net122)
  );
  and_cell and33 (
    .a (net119),
    .b (net121),
    .out (net126)
  );
  dffsr_cell flop15 (
    .d (net127),
    .clk (net1),
    .s (net128),
    .r (net104),
    .q (net129),
    .notq (net130)
  );
  mux_cell mux15 (
    .a (net129),
    .b (net130),
    .sel (net131),
    .out (net127)
  );
  and_cell and34 (
    .a (net124),
    .b (net126),
    .out (net131)
  );
  not_cell not1 (
    .in (net2),
    .out (net132)
  );
  dffsr_cell flop16 (
    .d (net133),
    .clk (net1),
    .s (net134),
    .r (net104),
    .q (net135),
    .notq (net136)
  );
  mux_cell mux16 (
    .a (net135),
    .b (net136),
    .sel (net137),
    .out (net133)
  );
  dffsr_cell flop17 (
    .d (net138),
    .clk (net1),
    .s (net139),
    .r (net104),
    .q (net140),
    .notq (net141)
  );
  mux_cell mux17 (
    .a (net140),
    .b (net141),
    .sel (net142),
    .out (net138)
  );
  and_cell and35 (
    .a (net135),
    .b (net137),
    .out (net142)
  );
  dffsr_cell flop18 (
    .d (net143),
    .clk (net1),
    .s (net144),
    .r (net104),
    .q (net145),
    .notq (net146)
  );
  mux_cell mux18 (
    .a (net145),
    .b (net146),
    .sel (net147),
    .out (net143)
  );
  and_cell and36 (
    .a (net140),
    .b (net142),
    .out (net147)
  );
  dffsr_cell flop19 (
    .d (net148),
    .clk (net1),
    .s (net149),
    .r (net104),
    .q (net150),
    .notq (net151)
  );
  mux_cell mux19 (
    .a (net150),
    .b (net151),
    .sel (net152),
    .out (net148)
  );
  and_cell and37 (
    .a (net145),
    .b (net147),
    .out (net152)
  );
  dffsr_cell flop20 (
    .d (net153),
    .clk (net1),
    .s (net154),
    .r (net104),
    .q (net155),
    .notq (net156)
  );
  mux_cell mux20 (
    .a (net155),
    .b (net156),
    .sel (net157),
    .out (net153)
  );
  and_cell and38 (
    .a (net150),
    .b (net152),
    .out (net157)
  );
  and_cell and39 (
    .a (net129),
    .b (net131),
    .out (net137)
  );
  dffsr_cell flop21 (
    .d (net158),
    .clk (net1),
    .s (net159),
    .r (net104),
    .q (net160),
    .notq (net161)
  );
  mux_cell mux21 (
    .a (net160),
    .b (net161),
    .sel (net162),
    .out (net158)
  );
  and_cell and40 (
    .a (net155),
    .b (net157),
    .out (net162)
  );
  dffsr_cell flop22 (
    .d (net163),
    .clk (net1),
    .s (net164),
    .r (net104),
    .q (net165),
    .notq (net166)
  );
  mux_cell mux22 (
    .a (net165),
    .b (net166),
    .sel (net167),
    .out (net163)
  );
  and_cell and41 (
    .a (net160),
    .b (net162),
    .out (net167)
  );
  dffsr_cell flop23 (
    .d (net168),
    .clk (net1),
    .s (net169),
    .r (net104),
    .q (net170),
    .notq (net171)
  );
  mux_cell mux23 (
    .a (net170),
    .b (net171),
    .sel (net172),
    .out (net168)
  );
  and_cell and42 (
    .a (net165),
    .b (net167),
    .out (net172)
  );
  dffsr_cell flop24 (
    .d (net173),
    .clk (net1),
    .s (net174),
    .r (net104),
    .q (net175),
    .notq (net176)
  );
  mux_cell mux24 (
    .a (net175),
    .b (net176),
    .sel (net177),
    .out (net173)
  );
  and_cell and43 (
    .a (net170),
    .b (net172),
    .out (net177)
  );
  dffsr_cell flop25 (
    .d (net178),
    .clk (net1),
    .s (net179),
    .r (net25),
    .q (net180),
    .notq ()
  );
  dffsr_cell flop26 (
    .d (net180),
    .clk (net1),
    .s (net179),
    .r (net25),
    .q (net181),
    .notq ()
  );
  dffsr_cell flop27 (
    .d (net181),
    .clk (net1),
    .s (net179),
    .r (net25),
    .q (),
    .notq (net182)
  );
  and_cell and64 (
    .a (net181),
    .b (net182),
    .out (net183)
  );
  xor_cell xor1 (
    .a (net10),
    .b (net175),
    .out (net184)
  );
  xor_cell xor2 (
    .a (net9),
    .b (net170),
    .out (net185)
  );
  xor_cell xor3 (
    .a (net8),
    .b (net165),
    .out (net186)
  );
  xor_cell xor4 (
    .a (net7),
    .b (net160),
    .out (net187)
  );
  xor_cell xor5 (
    .a (net6),
    .b (net155),
    .out (net188)
  );
  xor_cell xor6 (
    .a (net5),
    .b (net150),
    .out (net189)
  );
  xor_cell xor7 (
    .a (net4),
    .b (net145),
    .out (net190)
  );
  xor_cell xor8 (
    .a (net3),
    .b (net140),
    .out (net191)
  );
  and_cell and44 (
    .a (net192),
    .b (net193),
    .out (net194)
  );
  and_cell and45 (
    .a (net195),
    .b (net196),
    .out (net197)
  );
  and_cell and46 (
    .a (net198),
    .b (net199),
    .out (net200)
  );
  and_cell and47 (
    .a (net201),
    .b (net202),
    .out (net203)
  );
  and_cell and48 (
    .a (net200),
    .b (net203),
    .out (net204)
  );
  and_cell and49 (
    .a (net205),
    .b (net197),
    .out (net206)
  );
  and_cell and50 (
    .a (net206),
    .b (net204),
    .out (net178)
  );
  or_cell or1 (
    .a (net132),
    .b (net183),
    .out (net104)
  );
  not_cell not2 (
    .in (net184),
    .out (net202)
  );
  not_cell not3 (
    .in (net185),
    .out (net201)
  );
  not_cell not4 (
    .in (net187),
    .out (net198)
  );
  not_cell not6 (
    .in (net186),
    .out (net199)
  );
  not_cell not7 (
    .in (net189),
    .out (net195)
  );
  not_cell not8 (
    .in (net188),
    .out (net196)
  );
  not_cell not9 (
    .in (net191),
    .out (net192)
  );
  not_cell not10 (
    .in (net190),
    .out (net193)
  );
  dffsr_cell flop29 (
    .d (net207),
    .clk (net1),
    .s (net208),
    .r (net25),
    .q (net209),
    .notq (net210)
  );
  mux_cell mux25 (
    .a (net209),
    .b (net211),
    .sel (net45),
    .out (net207)
  );
  dffsr_cell flop30 (
    .d (net212),
    .clk (net1),
    .s (net213),
    .r (net25),
    .q (net214),
    .notq (net215)
  );
  dffsr_cell flop31 (
    .d (net216),
    .clk (net1),
    .s (net25),
    .r (net25),
    .q (net217),
    .notq ()
  );
  dffsr_cell flop32 (
    .d (net218),
    .clk (net1),
    .s (net213),
    .r (net25),
    .q (net219),
    .notq ()
  );
  dffsr_cell flop33 (
    .d (net220),
    .clk (net1),
    .s (net213),
    .r (net25),
    .q (net221),
    .notq ()
  );
  dffsr_cell flop34 (
    .d (net222),
    .clk (net1),
    .s (net213),
    .r (net25),
    .q (net223),
    .notq ()
  );
  dffsr_cell flop35 (
    .d (net224),
    .clk (net1),
    .s (net25),
    .r (net225),
    .q (net226),
    .notq ()
  );
  dffsr_cell flop36 (
    .d (net227),
    .clk (net1),
    .s (net213),
    .r (net25),
    .q (net228),
    .notq ()
  );
  dffsr_cell flop37 (
    .d (net229),
    .clk (net1),
    .s (net25),
    .r (net230),
    .q (net231),
    .notq ()
  );
  xor_cell xor11 (
    .a (net221),
    .b (net232),
    .out (net233)
  );
  and_cell and51 (
    .a (net210),
    .b (net59),
    .out (net234)
  );
  and_cell and52 (
    .a (net210),
    .b (net60),
    .out (net235)
  );
  and_cell and53 (
    .a (net210),
    .b (net62),
    .out (net236)
  );
  and_cell and54 (
    .a (net210),
    .b (net63),
    .out (net237)
  );
  and_cell and55 (
    .a (net210),
    .b (net65),
    .out (net238)
  );
  and_cell and56 (
    .a (net210),
    .b (net66),
    .out ()
  );
  and_cell and57 (
    .a (net210),
    .b (net67),
    .out (net239)
  );
  and_cell and58 (
    .a (net209),
    .b (net59),
    .out (net240)
  );
  and_cell and59 (
    .a (net209),
    .b (net60),
    .out (net241)
  );
  and_cell and60 (
    .a (net209),
    .b (net62),
    .out (net242)
  );
  and_cell and61 (
    .a (net209),
    .b (net63),
    .out (net243)
  );
  and_cell and62 (
    .a (net209),
    .b (net65),
    .out (net244)
  );
  and_cell and63 (
    .a (net209),
    .b (net66),
    .out (net245)
  );
  and_cell and65 (
    .a (net209),
    .b (net67),
    .out (net246)
  );
  or_cell or16 (
    .a (net236),
    .b (net234),
    .out (net247)
  );
  or_cell or17 (
    .a (net248),
    .b (net249),
    .out (net250)
  );
  and_cell and66 (
    .a (net235),
    .b (net214),
    .out (net249)
  );
  and_cell and67 (
    .a (net215),
    .b (net235),
    .out (net248)
  );
  or_cell or19 (
    .a (net237),
    .b (net248),
    .out (net251)
  );
  or_cell or20 (
    .a (net252),
    .b (net236),
    .out (net253)
  );
  and_cell and68 (
    .a (net238),
    .b (net214),
    .out (net252)
  );
  and_cell and69 (
    .a (net215),
    .b (net238),
    .out (net254)
  );
  or_cell or18 (
    .a (net254),
    .b (net252),
    .out (net255)
  );
  or_cell or21 (
    .a (net254),
    .b (net256),
    .out (net257)
  );
  and_cell and70 (
    .a (net239),
    .b (net214),
    .out (net258)
  );
  and_cell and71 (
    .a (net215),
    .b (net239),
    .out (net256)
  );
  or_cell or24 (
    .a (net259),
    .b (net240),
    .out (net260)
  );
  or_cell or25 (
    .a (net261),
    .b (net240),
    .out (net262)
  );
  or_cell or26 (
    .a (net243),
    .b (net261),
    .out (net263)
  );
  or_cell or27 (
    .a (net251),
    .b (net245),
    .out (net264)
  );
  and_cell and72 (
    .a (net242),
    .b (net214),
    .out (net265)
  );
  and_cell and73 (
    .a (net215),
    .b (net242),
    .out (net261)
  );
  or_cell or28 (
    .a (net244),
    .b (net265),
    .out (net266)
  );
  or_cell or29 (
    .a (net244),
    .b (net267),
    .out (net268)
  );
  and_cell and74 (
    .a (net245),
    .b (net214),
    .out (net267)
  );
  and_cell and75 (
    .a (net246),
    .b (net214),
    .out (net259)
  );
  and_cell and76 (
    .a (net215),
    .b (net246),
    .out (net269)
  );
  or_cell or31 (
    .a (net269),
    .b (net268),
    .out (net270)
  );
  or_cell or32 (
    .a (net256),
    .b (net258),
    .out (net271)
  );
  or_cell or22 (
    .a (net253),
    .b (net250),
    .out (net272)
  );
  or_cell or30 (
    .a (net266),
    .b (net260),
    .out (net273)
  );
  or_cell or33 (
    .a (net257),
    .b (net247),
    .out (net274)
  );
  or_cell or34 (
    .a (net273),
    .b (net274),
    .out (net275)
  );
  or_cell or35 (
    .a (net263),
    .b (net272),
    .out (net276)
  );
  or_cell or36 (
    .a (net270),
    .b (net276),
    .out (net277)
  );
  or_cell or37 (
    .a (net271),
    .b (net262),
    .out (net278)
  );
  or_cell or38 (
    .a (net255),
    .b (net264),
    .out (net279)
  );
  or_cell or39 (
    .a (net278),
    .b (net279),
    .out (net280)
  );
  dff_cell flop28 (
    .d (net95),
    .clk (net1),
    .q (net11),
    .notq ()
  );
  dff_cell flop46 (
    .d (net96),
    .clk (net1),
    .q (net12),
    .notq ()
  );
  dff_cell flop47 (
    .d (net97),
    .clk (net1),
    .q (net13),
    .notq ()
  );
  dff_cell flop48 (
    .d (net98),
    .clk (net1),
    .q (net14),
    .notq ()
  );
  dff_cell flop49 (
    .d (net99),
    .clk (net1),
    .q (net15),
    .notq ()
  );
  dff_cell flop50 (
    .d (net100),
    .clk (net1),
    .q (net16),
    .notq ()
  );
  dff_cell flop51 (
    .d (net101),
    .clk (net1),
    .q (net17),
    .notq ()
  );
  dff_cell flop52 (
    .d (net183),
    .clk (net1),
    .q (net45),
    .notq ()
  );
  dff_cell flop53 (
    .d (net275),
    .clk (net1),
    .q (net44),
    .notq ()
  );
  dff_cell flop54 (
    .d (net277),
    .clk (net1),
    .q (net46),
    .notq ()
  );
  dff_cell flop55 (
    .d (net280),
    .clk (net1),
    .q (net47),
    .notq ()
  );
  dff_cell flop56 (
    .d (net281),
    .clk (net1),
    .q (net211),
    .notq ()
  );
  mux_cell mux26 (
    .a (net214),
    .b (net233),
    .sel (net45),
    .out (net212)
  );
  mux_cell mux27 (
    .a (net217),
    .b (net214),
    .sel (net45),
    .out (net216)
  );
  mux_cell mux28 (
    .a (net219),
    .b (net217),
    .sel (net45),
    .out (net218)
  );
  mux_cell mux29 (
    .a (net221),
    .b (net219),
    .sel (net45),
    .out (net220)
  );
  mux_cell mux30 (
    .a (net223),
    .b (net221),
    .sel (net45),
    .out (net222)
  );
  xor_cell xor9 (
    .a (net223),
    .b (net282),
    .out (net232)
  );
  mux_cell mux31 (
    .a (net226),
    .b (net223),
    .sel (net45),
    .out (net224)
  );
  xor_cell xor10 (
    .a (net226),
    .b (net231),
    .out (net282)
  );
  mux_cell mux32 (
    .a (net228),
    .b (net226),
    .sel (net45),
    .out (net227)
  );
  mux_cell mux33 (
    .a (net231),
    .b (net228),
    .sel (net45),
    .out (net229)
  );
  or_cell or40 (
    .a (net240),
    .b (net241),
    .out (net283)
  );
  or_cell or41 (
    .a (net243),
    .b (net244),
    .out (net284)
  );
  or_cell or42 (
    .a (net283),
    .b (net284),
    .out (net285)
  );
  or_cell or43 (
    .a (net259),
    .b (net258),
    .out (net286)
  );
  or_cell or23 (
    .a (net285),
    .b (net286),
    .out (net287)
  );
  or_cell or44 (
    .a (net265),
    .b (net252),
    .out (net288)
  );
  or_cell or45 (
    .a (net287),
    .b (net289),
    .out (net281)
  );
  or_cell or46 (
    .a (net245),
    .b (net288),
    .out (net289)
  );
  and_cell and77 (
    .a (net135),
    .b (net194),
    .out (net205)
  );
endmodule
