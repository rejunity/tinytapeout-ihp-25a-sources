magic
tech sky130A
timestamp 1738436132
<< locali >>
rect -50 150000 50 150028
rect -50 -150028 50 -150000
<< rlocali >>
rect -50 -150000 50 150000
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 1.0 l 3000.0 m 1 nx 1 wmin 0.17 lmin 0.17 class resistor rho 12.8 val 38.4k dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
