magic
tech sky130A
magscale 1 2
timestamp 1738436334
<< error_p >>
rect 14571 646 14589 680
rect 14869 646 14904 680
rect 14571 -15 14588 646
rect 14870 627 14904 646
rect 14700 578 14758 584
rect 14700 544 14712 578
rect 14700 538 14758 544
rect 14700 68 14758 74
rect 14700 34 14712 68
rect 14700 28 14758 34
rect 14889 -68 14904 627
rect 14923 593 14958 627
rect 14923 -68 14957 593
rect 15069 525 15127 531
rect 15069 491 15081 525
rect 15069 485 15127 491
rect 15069 15 15127 21
rect 15069 -19 15081 15
rect 15069 -25 15127 -19
rect 14923 -102 14938 -68
<< error_s >>
rect 13682 1623 13717 1657
rect 13683 1604 13717 1623
rect 13491 1555 13553 1561
rect 13491 1521 13503 1555
rect 13491 1515 13553 1521
rect 13491 227 13553 233
rect 13491 193 13503 227
rect 13491 187 13553 193
rect 13702 91 13717 1604
rect 13736 1570 13771 1604
rect 14091 1570 14126 1604
rect 13736 91 13770 1570
rect 14092 1551 14126 1570
rect 13900 1502 13962 1508
rect 13900 1468 13912 1502
rect 13900 1462 13962 1468
rect 13900 174 13962 180
rect 13900 140 13912 174
rect 13900 134 13962 140
rect 13736 57 13751 91
rect 14111 38 14126 1551
rect 14145 1517 14180 1551
rect 14145 38 14179 1517
rect 14309 1449 14371 1455
rect 14309 1415 14321 1449
rect 14309 1409 14371 1415
rect 14501 716 14535 734
rect 14501 680 14551 716
rect 14309 121 14371 127
rect 14309 87 14321 121
rect 14309 81 14371 87
rect 14145 4 14160 38
rect 14518 -51 14551 680
<< error_ps >>
rect 14551 -51 14571 716
use sky130_fd_pr__res_generic_l1_QHFG3U  R1
timestamp 1738436132
transform 1 0 6819 0 1 299847
box -100 -300057 100 300057
use schmitt_trigger_ro  x1
timestamp 1738436067
transform 1 0 13250 0 1 636
box 41 -846 2428 1057
use sky130_fd_pr__cap_mim_m3_1_AHUHXA  XC1
timestamp 1738436132
transform 1 0 10105 0 1 2830
box -3186 -3040 3186 3040
<< end >>
