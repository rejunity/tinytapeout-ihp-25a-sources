magic
tech sky130A
magscale 1 2
timestamp 1738434555
<< checkpaint >>
rect -1313 1358 2547 1646
rect -1313 1305 4252 1358
rect -1313 1252 4661 1305
rect -1313 1199 5070 1252
rect -1313 1146 5479 1199
rect -1313 987 5888 1146
rect -1313 828 7035 987
rect -1313 -1843 8182 828
rect -1313 -2214 2547 -1843
rect 2906 -1896 8182 -1843
rect 4053 -2055 8182 -1896
rect 5200 -2214 8182 -2055
<< error_s >>
rect 298 381 333 415
rect 299 362 333 381
rect 129 313 187 319
rect 129 279 141 313
rect 129 273 187 279
rect 129 119 187 125
rect 129 85 141 119
rect 129 79 187 85
rect 318 -17 333 362
rect 352 328 387 362
rect 667 328 702 362
rect 352 -17 386 328
rect 668 309 702 328
rect 498 260 556 266
rect 498 226 510 260
rect 498 220 556 226
rect 498 66 556 72
rect 498 32 510 66
rect 498 26 556 32
rect 352 -51 367 -17
rect 687 -70 702 309
rect 721 275 756 309
rect 1036 275 1071 309
rect 721 -70 755 275
rect 1037 256 1071 275
rect 867 207 925 213
rect 867 173 879 207
rect 867 167 925 173
rect 867 13 925 19
rect 867 -21 879 13
rect 867 -27 925 -21
rect 721 -104 736 -70
rect 1056 -123 1071 256
rect 1090 222 1125 256
rect 1405 222 1440 256
rect 1090 -123 1124 222
rect 1406 203 1440 222
rect 1236 154 1294 160
rect 1236 120 1248 154
rect 1236 114 1294 120
rect 1236 -40 1294 -34
rect 1236 -74 1248 -40
rect 1236 -80 1294 -74
rect 1090 -157 1105 -123
rect 1425 -176 1440 203
rect 1459 169 1494 203
rect 1774 169 1809 203
rect 1459 -176 1493 169
rect 1775 150 1809 169
rect 1605 101 1663 107
rect 1605 67 1617 101
rect 1605 61 1663 67
rect 1605 -93 1663 -87
rect 1605 -127 1617 -93
rect 1605 -133 1663 -127
rect 1459 -210 1474 -176
rect 1794 -229 1809 150
rect 1828 116 1863 150
rect 2143 116 2178 150
rect 1828 -229 1862 116
rect 2144 97 2178 116
rect 2530 97 2583 98
rect 1974 48 2032 54
rect 1974 14 1986 48
rect 1974 8 2032 14
rect 1974 -146 2032 -140
rect 1974 -180 1986 -146
rect 1974 -186 2032 -180
rect 1828 -263 1843 -229
rect 2163 -282 2178 97
rect 2197 63 2232 97
rect 2512 63 2583 97
rect 2197 -282 2231 63
rect 2513 62 2583 63
rect 2530 28 2601 62
rect 2921 28 2956 62
rect 2343 -5 2401 1
rect 2343 -39 2355 -5
rect 2343 -45 2401 -39
rect 2343 -199 2401 -193
rect 2343 -233 2355 -199
rect 2343 -239 2401 -233
rect 2197 -316 2212 -282
rect 2530 -335 2600 28
rect 2922 9 2956 28
rect 2730 -40 2792 -34
rect 2730 -74 2742 -40
rect 2730 -80 2792 -74
rect 2730 -252 2792 -246
rect 2730 -286 2742 -252
rect 2730 -292 2792 -286
rect 2530 -371 2583 -335
rect 2941 -388 2956 9
rect 2975 -25 3010 9
rect 3330 -25 3365 9
rect 2975 -388 3009 -25
rect 3331 -44 3365 -25
rect 3139 -93 3201 -87
rect 3139 -127 3151 -93
rect 3139 -133 3201 -127
rect 3139 -305 3201 -299
rect 3139 -339 3151 -305
rect 3139 -345 3201 -339
rect 2975 -422 2990 -388
rect 3350 -441 3365 -44
rect 3384 -78 3419 -44
rect 3739 -78 3774 -44
rect 3384 -441 3418 -78
rect 3740 -97 3774 -78
rect 3548 -146 3610 -140
rect 3548 -180 3560 -146
rect 3548 -186 3610 -180
rect 3548 -358 3610 -352
rect 3548 -392 3560 -358
rect 3548 -398 3610 -392
rect 3384 -475 3399 -441
rect 3759 -494 3774 -97
rect 3793 -131 3828 -97
rect 4148 -131 4183 -97
rect 3793 -494 3827 -131
rect 4149 -150 4183 -131
rect 3957 -199 4019 -193
rect 3957 -233 3969 -199
rect 3957 -239 4019 -233
rect 3957 -411 4019 -405
rect 3957 -445 3969 -411
rect 3957 -451 4019 -445
rect 3793 -528 3808 -494
rect 4168 -547 4183 -150
rect 4202 -184 4237 -150
rect 4557 -184 4592 -167
rect 4202 -547 4236 -184
rect 4558 -185 4592 -184
rect 4558 -221 4628 -185
rect 4366 -252 4428 -246
rect 4366 -286 4378 -252
rect 4575 -255 4646 -221
rect 4926 -255 4961 -221
rect 4366 -292 4428 -286
rect 4366 -464 4428 -458
rect 4366 -498 4378 -464
rect 4366 -504 4428 -498
rect 4202 -581 4217 -547
rect 4575 -600 4645 -255
rect 4927 -274 4961 -255
rect 5313 -274 5366 -273
rect 4757 -323 4815 -317
rect 4757 -357 4769 -323
rect 4757 -363 4815 -357
rect 4757 -517 4815 -511
rect 4757 -551 4769 -517
rect 4757 -557 4815 -551
rect 4575 -636 4628 -600
rect 4946 -653 4961 -274
rect 4980 -308 5015 -274
rect 5295 -308 5366 -274
rect 4980 -653 5014 -308
rect 5296 -309 5366 -308
rect 5313 -343 5384 -309
rect 5704 -343 5739 -326
rect 5126 -376 5184 -370
rect 5126 -410 5138 -376
rect 5126 -416 5184 -410
rect 5126 -570 5184 -564
rect 5126 -604 5138 -570
rect 5126 -610 5184 -604
rect 4980 -687 4995 -653
rect 5313 -706 5383 -343
rect 5705 -344 5739 -343
rect 5705 -380 5775 -344
rect 5513 -411 5575 -405
rect 5513 -445 5525 -411
rect 5722 -414 5793 -380
rect 6073 -414 6108 -380
rect 5513 -451 5575 -445
rect 5513 -623 5575 -617
rect 5513 -657 5525 -623
rect 5513 -663 5575 -657
rect 5313 -742 5366 -706
rect 5722 -759 5792 -414
rect 6074 -433 6108 -414
rect 5904 -482 5962 -476
rect 5904 -516 5916 -482
rect 5904 -522 5962 -516
rect 5904 -676 5962 -670
rect 5904 -710 5916 -676
rect 5904 -716 5962 -710
rect 5722 -795 5775 -759
rect 6093 -812 6108 -433
rect 6127 -467 6162 -433
rect 6127 -812 6161 -467
rect 6273 -535 6331 -529
rect 6273 -569 6285 -535
rect 6273 -575 6331 -569
rect 6273 -729 6331 -723
rect 6273 -763 6285 -729
rect 6273 -769 6331 -763
rect 6127 -846 6142 -812
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM1
timestamp 0
transform 1 0 158 0 1 199
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM2
timestamp 0
transform 1 0 527 0 1 146
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM3
timestamp 0
transform 1 0 896 0 1 93
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM4
timestamp 0
transform 1 0 1265 0 1 40
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM5
timestamp 0
transform 1 0 1634 0 1 -13
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM6
timestamp 0
transform 1 0 2003 0 1 -66
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XM7
timestamp 0
transform 1 0 2372 0 1 -119
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XM8
timestamp 0
transform 1 0 2761 0 1 -163
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XM9
timestamp 0
transform 1 0 3170 0 1 -216
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XM10
timestamp 0
transform 1 0 3579 0 1 -269
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XM11
timestamp 0
transform 1 0 3988 0 1 -322
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XM12
timestamp 0
transform 1 0 4397 0 1 -375
box -231 -261 231 261
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XMa
timestamp 0
transform 1 0 5544 0 1 -534
box -231 -261 231 261
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XMb
timestamp 0
transform 1 0 5155 0 1 -490
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XMc
timestamp 0
transform 1 0 4786 0 1 -437
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_lvt_A33RKA  XMd
timestamp 0
transform 1 0 6691 0 1 -693
box -231 -261 231 261
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XMe
timestamp 0
transform 1 0 6302 0 1 -649
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_lvt_BK97Z7  XMf
timestamp 0
transform 1 0 5933 0 1 -596
box -211 -252 211 252
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 -53 0 1 -954
box 0 0 1340 1340
<< end >>
