** sch_path: /foss/designs/tt10-uR-IPs/xschem/T3/oscillators/A_tt10_Ring_currentStarved/osc_general_tran_tb.sch
**.subckt osc_general_tran_tb
VIN1 net2 0 0 pulse 0 1.8 100u 1u 1u 1 2 ac 1 0
vi_total net1 Vjump 0
.save i(vi_total)
R2 net1 net2 30 m=1
C1 Vclk 0 1f m=1
x1 net9 net10 net6 Vclk net5 osc
vi_bias_n net7 0 0
.save i(vi_bias_n)
vi_bias_p Vjump net8 0
.save i(vi_bias_p)
vi_3 net3 net5 0
.save i(vi_3)
vi_4 net4 net6 0
.save i(vi_4)
vi_osc_p Vjump net9 0
.save i(vi_osc_p)
vi_osc_n 0 net10 0
.save i(vi_osc_n)
x2 net8 net7 net3 net4 ibias_10nA_parax
**** begin user architecture code



.temp 30
.param Vdd = 1.8
.param imax = 100e-9


.option savecurrents
.save all
.control
  save all alli
  save

  op
  write osc_51k5Hz_tb.raw
  remzerovec
  set appendwrite

  tran 0.1u 1.5m
  remzerovec
  write osc_51k5Hz_tb.raw





  *quit 0




.endc




** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  T3/oscillators/A_tt10_Ring_currentStarved/osc.sym # of pins=5
** sym_path: /foss/designs/tt10-uR-IPs/xschem/T3/oscillators/A_tt10_Ring_currentStarved/osc.sym
** sch_path: /foss/designs/tt10-uR-IPs/xschem/T3/oscillators/A_tt10_Ring_currentStarved/osc.sch
.subckt osc Vdd Vss pBias Out nBias
*.ipin Vdd
*.ipin Vss
*.opin Out
*.ipin nBias
*.ipin pBias
XM6 net1 nBias Vss Vss sky130_fd_pr__nfet_01v8 L=0.4 W=2.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net4 pBias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net2 nBias Vss Vss sky130_fd_pr__nfet_01v8 L=0.4 W=2.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net5 pBias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net3 nBias Vss Vss sky130_fd_pr__nfet_01v8 L=0.4 W=2.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net6 pBias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 net10 net2 net5 net11 Vdd Vss schmTrigg
x1 net7 net1 net4 net10 Vdd Vss schmTrigg
x4 net11 net3 net6 net7 Vdd Vss schmTrigg
XM1 net8 nBias Vss Vss sky130_fd_pr__nfet_01v8 L=0.4 W=2.25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net9 pBias Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x5 net7 net8 net9 Out Vdd Vss schmTrigg
XC1 net10 Vss sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XC2 net11 Vss sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XC3 net7 Vss sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  T2/biasGen/A_tt10_10nA/ibias_10nA_parax.sym # of pins=4
** sym_path: /foss/designs/tt10-uR-IPs/xschem/T2/biasGen/A_tt10_10nA/ibias_10nA_parax.sym
.include T2/biasGen/A_tt10_10nA/ibias_10nA_parax.spice

* expanding   symbol:  T1/schmTrigg/schmTrigg.sym # of pins=6
** sym_path: /foss/designs/tt10-uR-IPs/xschem/T1/schmTrigg/schmTrigg.sym
** sch_path: /foss/designs/tt10-uR-IPs/xschem/T1/schmTrigg/schmTrigg.sch
.subckt schmTrigg Vin VSS VDD Vout pBulk nBulk
*.ipin Vin
*.ipin VDD
*.ipin VSS
*.opin Vout
*.ipin nBulk
*.ipin pBulk
XM1 VDD Vout Vn nBulk sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vn Vin VSS nBulk sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout Vin Vn nBulk sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 VSS Vout Vp pBulk sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vout Vin Vp pBulk sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vp Vin VDD pBulk sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
