magic
tech sky130A
magscale 1 2
timestamp 1741535882
<< metal4 >>
rect -849 539 849 580
rect -849 -539 593 539
rect 829 -539 849 539
rect -849 -580 849 -539
<< via4 >>
rect 593 -539 829 539
<< mimcap2 >>
rect -769 460 231 500
rect -769 -460 -729 460
rect 191 -460 231 460
rect -769 -500 231 -460
<< mimcap2contact >>
rect -729 -460 191 460
<< metal5 >>
rect 551 539 871 581
rect -753 460 215 484
rect -753 -460 -729 460
rect 191 -460 215 460
rect -753 -484 215 -460
rect 551 -539 593 539
rect 829 -539 871 539
rect 551 -581 871 -539
<< properties >>
string FIXED_BBOX -849 -580 311 580
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 5 l 5 val 53.8 carea 2.00 cperi 0.19 class capacitor nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
