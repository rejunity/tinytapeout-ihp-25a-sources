`default_nettype none
module barrier_rom(
    input  wire [3:0] row_index,   
    output wire [31:0] row_data    
);
    reg [31:0] rom_array [0:15];
    initial begin
        // Example barrier pattern. Customize as needed.
        rom_array[0]  = 32'b00000111111111111111111111100000;
        rom_array[1]  = 32'b00001111111111111111111111110000;
        rom_array[2]  = 32'b00011111111111111111111111111000;
        rom_array[3]  = 32'b00111111111111111111111111111100;
        rom_array[4]  = 32'b01111111111111111111111111111110;
        rom_array[5]  = 32'b11111111111111111111111111111111;
        rom_array[6]  = 32'b11111111111111111111111111111111;
        rom_array[7]  = 32'b11111111111111111111111111111111;
        rom_array[8]  = 32'b11111111111111111111111111111111;
        rom_array[9]  = 32'b11111111111111111111111111111111;
        rom_array[10] = 32'b11111111111111111111111111111111;
        rom_array[11] = 32'b11111111111111111111111111111111;
        rom_array[12] = 32'b11111111111111111111111111111111;
        rom_array[13] = 32'b11111111100000000000000111111111;
        rom_array[14] = 32'b11111111000000000000000011111111;
        rom_array[15] = 32'b11111110000000000000000001111111;
    end
    assign row_data = rom_array[row_index];
endmodule