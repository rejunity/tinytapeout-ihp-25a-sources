/* Automatically generated from https://wokwi.com/projects/414118423095874561 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_414118423095874561(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = ui_in[0];
  wire net3;
  wire net4;
  wire net5 = 1'b0;
  wire net6 = 1'b1;
  wire net7 = 1'b1;
  wire net8 = 1'b0;
  wire net9 = 1'b1;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;
  wire net474;
  wire net475;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;

  assign uo_out[0] = 0;
  assign uo_out[1] = net3;
  assign uo_out[2] = net3;
  assign uo_out[3] = net3;
  assign uo_out[4] = net3;
  assign uo_out[5] = net3;
  assign uo_out[6] = 0;
  assign uo_out[7] = net4;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  dff_cell flop1 (
    .d (net2),
    .clk (net10),
    .q (net3),
    .notq (net11)
  );
  dff_cell flop2 (
    .d (net12),
    .clk (net10),
    .q (net13),
    .notq ()
  );
  dff_cell flop3 (
    .d (net14),
    .clk (net1),
    .q (net15),
    .notq ()
  );
  dff_cell flop4 (
    .d (net13),
    .clk (net1),
    .q (net14),
    .notq ()
  );
  dff_cell flop5 (
    .d (net15),
    .clk (net1),
    .q (net16),
    .notq ()
  );
  dff_cell flop6 (
    .d (net17),
    .clk (net1),
    .q (net18),
    .notq ()
  );
  dff_cell flop7 (
    .d (net19),
    .clk (net20),
    .q (net21),
    .notq ()
  );
  dff_cell flop8 (
    .d (net22),
    .clk (net18),
    .q (net23),
    .notq (net20)
  );
  dff_cell flop9 (
    .d (net24),
    .clk (net21),
    .q (net25),
    .notq ()
  );
  not_cell not1 (
    .in (net18),
    .out (net17)
  );
  not_cell not2 (
    .in (net23),
    .out (net22)
  );
  not_cell not3 (
    .in (net21),
    .out (net19)
  );
  not_cell not4 (
    .in (net25),
    .out (net24)
  );
  dff_cell flop10 (
    .d (net26),
    .clk (net25),
    .q (net27),
    .notq ()
  );
  dff_cell flop11 (
    .d (net28),
    .clk (net29),
    .q (net30),
    .notq ()
  );
  dff_cell flop12 (
    .d (net31),
    .clk (net27),
    .q (net32),
    .notq (net29)
  );
  dff_cell flop13 (
    .d (net33),
    .clk (net30),
    .q (net34),
    .notq ()
  );
  not_cell not5 (
    .in (net27),
    .out (net26)
  );
  not_cell not6 (
    .in (net32),
    .out (net31)
  );
  not_cell not7 (
    .in (net30),
    .out (net28)
  );
  not_cell not8 (
    .in (net34),
    .out (net33)
  );
  dff_cell flop14 (
    .d (net35),
    .clk (net34),
    .q (net36),
    .notq ()
  );
  dff_cell flop15 (
    .d (net37),
    .clk (net38),
    .q (net39),
    .notq ()
  );
  dff_cell flop16 (
    .d (net40),
    .clk (net36),
    .q (net41),
    .notq (net38)
  );
  dff_cell flop17 (
    .d (net42),
    .clk (net39),
    .q (net43),
    .notq ()
  );
  not_cell not9 (
    .in (net36),
    .out (net35)
  );
  not_cell not10 (
    .in (net41),
    .out (net40)
  );
  not_cell not11 (
    .in (net39),
    .out (net37)
  );
  not_cell not12 (
    .in (net43),
    .out (net42)
  );
  dff_cell flop18 (
    .d (net44),
    .clk (net43),
    .q (net45),
    .notq ()
  );
  dff_cell flop19 (
    .d (net46),
    .clk (net47),
    .q (net48),
    .notq ()
  );
  dff_cell flop20 (
    .d (net49),
    .clk (net45),
    .q (net50),
    .notq (net47)
  );
  dff_cell flop21 (
    .d (net51),
    .clk (net48),
    .q (net52),
    .notq ()
  );
  not_cell not13 (
    .in (net45),
    .out (net44)
  );
  not_cell not14 (
    .in (net50),
    .out (net49)
  );
  not_cell not15 (
    .in (net48),
    .out (net46)
  );
  not_cell not16 (
    .in (net52),
    .out (net51)
  );
  dff_cell flop22 (
    .d (net53),
    .clk (net52),
    .q (net54),
    .notq ()
  );
  dff_cell flop23 (
    .d (net55),
    .clk (net56),
    .q (net57),
    .notq ()
  );
  dff_cell flop24 (
    .d (net58),
    .clk (net54),
    .q (net59),
    .notq (net56)
  );
  dff_cell flop25 (
    .d (net60),
    .clk (net57),
    .q (net61),
    .notq ()
  );
  not_cell not17 (
    .in (net54),
    .out (net53)
  );
  not_cell not18 (
    .in (net59),
    .out (net58)
  );
  not_cell not19 (
    .in (net57),
    .out (net55)
  );
  not_cell not20 (
    .in (net61),
    .out (net60)
  );
  dff_cell flop26 (
    .d (net62),
    .clk (net61),
    .q (net63),
    .notq ()
  );
  dff_cell flop27 (
    .d (net64),
    .clk (net65),
    .q (net66),
    .notq ()
  );
  dff_cell flop28 (
    .d (net67),
    .clk (net63),
    .q (net68),
    .notq (net65)
  );
  dff_cell flop29 (
    .d (net69),
    .clk (net66),
    .q (net70),
    .notq ()
  );
  not_cell not21 (
    .in (net63),
    .out (net62)
  );
  not_cell not22 (
    .in (net68),
    .out (net67)
  );
  not_cell not23 (
    .in (net66),
    .out (net64)
  );
  not_cell not24 (
    .in (net70),
    .out (net69)
  );
  dff_cell flop30 (
    .d (net71),
    .clk (net70),
    .q (net72),
    .notq ()
  );
  dff_cell flop31 (
    .d (net73),
    .clk (net74),
    .q (net75),
    .notq ()
  );
  dff_cell flop32 (
    .d (net76),
    .clk (net72),
    .q (net77),
    .notq (net74)
  );
  dff_cell flop33 (
    .d (net78),
    .clk (net75),
    .q (net79),
    .notq ()
  );
  not_cell not25 (
    .in (net72),
    .out (net71)
  );
  not_cell not26 (
    .in (net77),
    .out (net76)
  );
  not_cell not27 (
    .in (net75),
    .out (net73)
  );
  not_cell not28 (
    .in (net79),
    .out (net78)
  );
  dff_cell flop34 (
    .d (net80),
    .clk (net79),
    .q (net81),
    .notq ()
  );
  dff_cell flop35 (
    .d (net82),
    .clk (net83),
    .q (net84),
    .notq ()
  );
  dff_cell flop36 (
    .d (net85),
    .clk (net81),
    .q (net86),
    .notq (net83)
  );
  dff_cell flop37 (
    .d (net87),
    .clk (net84),
    .q (net88),
    .notq ()
  );
  not_cell not29 (
    .in (net81),
    .out (net80)
  );
  not_cell not30 (
    .in (net86),
    .out (net85)
  );
  not_cell not31 (
    .in (net84),
    .out (net82)
  );
  not_cell not32 (
    .in (net88),
    .out (net87)
  );
  dff_cell flop38 (
    .d (net89),
    .clk (net88),
    .q (net90),
    .notq ()
  );
  dff_cell flop39 (
    .d (net91),
    .clk (net92),
    .q (net93),
    .notq ()
  );
  dff_cell flop40 (
    .d (net94),
    .clk (net90),
    .q (net95),
    .notq (net92)
  );
  dff_cell flop41 (
    .d (net96),
    .clk (net93),
    .q (net10),
    .notq ()
  );
  not_cell not33 (
    .in (net90),
    .out (net89)
  );
  not_cell not34 (
    .in (net95),
    .out (net94)
  );
  not_cell not35 (
    .in (net93),
    .out (net91)
  );
  not_cell not36 (
    .in (net10),
    .out (net96)
  );
  not_cell not37 (
    .in (net16),
    .out (net12)
  );
  not_cell not38 (
    .in (net97),
    .out (net98)
  );
  not_cell not39 (
    .in (net98),
    .out (net99)
  );
  not_cell not40 (
    .in (net99),
    .out (net100)
  );
  not_cell not41 (
    .in (net100),
    .out (net101)
  );
  not_cell not42 (
    .in (net102),
    .out (net103)
  );
  not_cell not43 (
    .in (net103),
    .out (net104)
  );
  not_cell not44 (
    .in (net104),
    .out (net105)
  );
  not_cell not45 (
    .in (net105),
    .out (net97)
  );
  not_cell not46 (
    .in (net106),
    .out (net107)
  );
  not_cell not47 (
    .in (net107),
    .out (net108)
  );
  not_cell not48 (
    .in (net108),
    .out (net109)
  );
  not_cell not49 (
    .in (net109),
    .out (net110)
  );
  not_cell not50 (
    .in (net101),
    .out (net111)
  );
  not_cell not51 (
    .in (net111),
    .out (net112)
  );
  not_cell not52 (
    .in (net112),
    .out (net113)
  );
  not_cell not53 (
    .in (net113),
    .out (net106)
  );
  not_cell not54 (
    .in (net114),
    .out (net115)
  );
  not_cell not55 (
    .in (net115),
    .out (net116)
  );
  not_cell not56 (
    .in (net116),
    .out (net117)
  );
  not_cell not57 (
    .in (net117),
    .out (net118)
  );
  not_cell not58 (
    .in (net110),
    .out (net119)
  );
  not_cell not59 (
    .in (net119),
    .out (net120)
  );
  not_cell not60 (
    .in (net120),
    .out (net121)
  );
  not_cell not61 (
    .in (net121),
    .out (net114)
  );
  not_cell not62 (
    .in (net122),
    .out (net123)
  );
  not_cell not63 (
    .in (net123),
    .out (net124)
  );
  not_cell not64 (
    .in (net124),
    .out (net125)
  );
  not_cell not65 (
    .in (net125),
    .out (net126)
  );
  not_cell not66 (
    .in (net118),
    .out (net127)
  );
  not_cell not67 (
    .in (net127),
    .out (net128)
  );
  not_cell not68 (
    .in (net128),
    .out (net129)
  );
  not_cell not69 (
    .in (net129),
    .out (net122)
  );
  not_cell not70 (
    .in (net130),
    .out (net131)
  );
  not_cell not71 (
    .in (net131),
    .out (net132)
  );
  not_cell not72 (
    .in (net132),
    .out (net133)
  );
  not_cell not73 (
    .in (net133),
    .out (net134)
  );
  not_cell not74 (
    .in (net80),
    .out (net135)
  );
  not_cell not75 (
    .in (net135),
    .out (net136)
  );
  not_cell not76 (
    .in (net136),
    .out (net137)
  );
  not_cell not77 (
    .in (net137),
    .out (net130)
  );
  not_cell not78 (
    .in (net138),
    .out (net139)
  );
  not_cell not79 (
    .in (net139),
    .out (net140)
  );
  not_cell not80 (
    .in (net140),
    .out (net141)
  );
  not_cell not81 (
    .in (net141),
    .out (net142)
  );
  not_cell not82 (
    .in (net134),
    .out (net143)
  );
  not_cell not83 (
    .in (net143),
    .out (net144)
  );
  not_cell not84 (
    .in (net144),
    .out (net145)
  );
  not_cell not85 (
    .in (net145),
    .out (net138)
  );
  not_cell not86 (
    .in (net146),
    .out (net147)
  );
  not_cell not87 (
    .in (net147),
    .out (net148)
  );
  not_cell not88 (
    .in (net148),
    .out (net149)
  );
  not_cell not89 (
    .in (net149),
    .out (net150)
  );
  not_cell not90 (
    .in (net142),
    .out (net151)
  );
  not_cell not91 (
    .in (net151),
    .out (net152)
  );
  not_cell not92 (
    .in (net152),
    .out (net153)
  );
  not_cell not93 (
    .in (net153),
    .out (net146)
  );
  not_cell not94 (
    .in (net154),
    .out (net155)
  );
  not_cell not95 (
    .in (net155),
    .out (net156)
  );
  not_cell not96 (
    .in (net156),
    .out (net157)
  );
  not_cell not97 (
    .in (net157),
    .out (net102)
  );
  not_cell not98 (
    .in (net150),
    .out (net158)
  );
  not_cell not99 (
    .in (net158),
    .out (net159)
  );
  not_cell not100 (
    .in (net159),
    .out (net160)
  );
  not_cell not101 (
    .in (net160),
    .out (net154)
  );
  not_cell not102 (
    .in (net161),
    .out (net162)
  );
  not_cell not103 (
    .in (net162),
    .out (net163)
  );
  not_cell not104 (
    .in (net163),
    .out (net164)
  );
  not_cell not105 (
    .in (net164),
    .out (net165)
  );
  not_cell not106 (
    .in (net166),
    .out (net167)
  );
  not_cell not107 (
    .in (net167),
    .out (net168)
  );
  not_cell not108 (
    .in (net168),
    .out (net169)
  );
  not_cell not109 (
    .in (net169),
    .out (net161)
  );
  not_cell not110 (
    .in (net170),
    .out (net171)
  );
  not_cell not111 (
    .in (net171),
    .out (net172)
  );
  not_cell not112 (
    .in (net172),
    .out (net173)
  );
  not_cell not113 (
    .in (net173),
    .out (net174)
  );
  not_cell not114 (
    .in (net165),
    .out (net175)
  );
  not_cell not115 (
    .in (net175),
    .out (net176)
  );
  not_cell not116 (
    .in (net176),
    .out (net177)
  );
  not_cell not117 (
    .in (net177),
    .out (net170)
  );
  not_cell not118 (
    .in (net178),
    .out (net179)
  );
  not_cell not119 (
    .in (net179),
    .out (net180)
  );
  not_cell not120 (
    .in (net180),
    .out (net181)
  );
  not_cell not121 (
    .in (net181),
    .out (net182)
  );
  not_cell not122 (
    .in (net174),
    .out (net183)
  );
  not_cell not123 (
    .in (net183),
    .out (net184)
  );
  not_cell not124 (
    .in (net184),
    .out (net185)
  );
  not_cell not125 (
    .in (net185),
    .out (net178)
  );
  not_cell not126 (
    .in (net186),
    .out (net187)
  );
  not_cell not127 (
    .in (net187),
    .out (net188)
  );
  not_cell not128 (
    .in (net188),
    .out (net189)
  );
  not_cell not129 (
    .in (net189),
    .out (net190)
  );
  not_cell not130 (
    .in (net182),
    .out (net191)
  );
  not_cell not131 (
    .in (net191),
    .out (net192)
  );
  not_cell not132 (
    .in (net192),
    .out (net193)
  );
  not_cell not133 (
    .in (net193),
    .out (net186)
  );
  not_cell not134 (
    .in (net194),
    .out (net195)
  );
  not_cell not135 (
    .in (net195),
    .out (net196)
  );
  not_cell not136 (
    .in (net196),
    .out (net197)
  );
  not_cell not137 (
    .in (net197),
    .out (net198)
  );
  not_cell not138 (
    .in (net126),
    .out (net199)
  );
  not_cell not139 (
    .in (net199),
    .out (net200)
  );
  not_cell not140 (
    .in (net200),
    .out (net201)
  );
  not_cell not141 (
    .in (net201),
    .out (net194)
  );
  not_cell not142 (
    .in (net202),
    .out (net203)
  );
  not_cell not143 (
    .in (net203),
    .out (net204)
  );
  not_cell not144 (
    .in (net204),
    .out (net205)
  );
  not_cell not145 (
    .in (net205),
    .out (net206)
  );
  not_cell not146 (
    .in (net198),
    .out (net207)
  );
  not_cell not147 (
    .in (net207),
    .out (net208)
  );
  not_cell not148 (
    .in (net208),
    .out (net209)
  );
  not_cell not149 (
    .in (net209),
    .out (net202)
  );
  not_cell not150 (
    .in (net210),
    .out (net211)
  );
  not_cell not151 (
    .in (net211),
    .out (net212)
  );
  not_cell not152 (
    .in (net212),
    .out (net213)
  );
  not_cell not153 (
    .in (net213),
    .out (net214)
  );
  not_cell not154 (
    .in (net206),
    .out (net215)
  );
  not_cell not155 (
    .in (net215),
    .out (net216)
  );
  not_cell not156 (
    .in (net216),
    .out (net217)
  );
  not_cell not157 (
    .in (net217),
    .out (net210)
  );
  not_cell not158 (
    .in (net218),
    .out (net219)
  );
  not_cell not159 (
    .in (net219),
    .out (net220)
  );
  not_cell not160 (
    .in (net220),
    .out (net221)
  );
  not_cell not161 (
    .in (net221),
    .out (net166)
  );
  not_cell not162 (
    .in (net214),
    .out (net222)
  );
  not_cell not163 (
    .in (net222),
    .out (net223)
  );
  not_cell not164 (
    .in (net223),
    .out (net224)
  );
  not_cell not165 (
    .in (net224),
    .out (net218)
  );
  not_cell not166 (
    .in (net225),
    .out (net226)
  );
  not_cell not167 (
    .in (net226),
    .out (net227)
  );
  not_cell not168 (
    .in (net227),
    .out (net228)
  );
  not_cell not169 (
    .in (net228),
    .out (net229)
  );
  not_cell not170 (
    .in (net230),
    .out (net231)
  );
  not_cell not171 (
    .in (net231),
    .out (net232)
  );
  not_cell not172 (
    .in (net232),
    .out (net233)
  );
  not_cell not173 (
    .in (net233),
    .out (net225)
  );
  not_cell not174 (
    .in (net234),
    .out (net235)
  );
  not_cell not175 (
    .in (net235),
    .out (net236)
  );
  not_cell not176 (
    .in (net236),
    .out (net237)
  );
  not_cell not177 (
    .in (net237),
    .out (net238)
  );
  not_cell not178 (
    .in (net229),
    .out (net239)
  );
  not_cell not179 (
    .in (net239),
    .out (net240)
  );
  not_cell not180 (
    .in (net240),
    .out (net241)
  );
  not_cell not181 (
    .in (net241),
    .out (net234)
  );
  not_cell not182 (
    .in (net242),
    .out (net243)
  );
  not_cell not183 (
    .in (net243),
    .out (net244)
  );
  not_cell not184 (
    .in (net244),
    .out (net245)
  );
  not_cell not185 (
    .in (net245),
    .out (net246)
  );
  not_cell not186 (
    .in (net238),
    .out (net247)
  );
  not_cell not187 (
    .in (net247),
    .out (net248)
  );
  not_cell not188 (
    .in (net248),
    .out (net249)
  );
  not_cell not189 (
    .in (net249),
    .out (net242)
  );
  not_cell not190 (
    .in (net250),
    .out (net251)
  );
  not_cell not191 (
    .in (net251),
    .out (net252)
  );
  not_cell not192 (
    .in (net252),
    .out (net253)
  );
  not_cell not193 (
    .in (net253),
    .out (net254)
  );
  not_cell not194 (
    .in (net246),
    .out (net255)
  );
  not_cell not195 (
    .in (net255),
    .out (net256)
  );
  not_cell not196 (
    .in (net256),
    .out (net257)
  );
  not_cell not197 (
    .in (net257),
    .out (net250)
  );
  not_cell not198 (
    .in (net258),
    .out (net259)
  );
  not_cell not199 (
    .in (net259),
    .out (net260)
  );
  not_cell not200 (
    .in (net260),
    .out (net261)
  );
  not_cell not201 (
    .in (net261),
    .out (net262)
  );
  not_cell not202 (
    .in (net190),
    .out (net263)
  );
  not_cell not203 (
    .in (net263),
    .out (net264)
  );
  not_cell not204 (
    .in (net264),
    .out (net265)
  );
  not_cell not205 (
    .in (net265),
    .out (net258)
  );
  not_cell not206 (
    .in (net266),
    .out (net267)
  );
  not_cell not207 (
    .in (net267),
    .out (net268)
  );
  not_cell not208 (
    .in (net268),
    .out (net269)
  );
  not_cell not209 (
    .in (net269),
    .out (net270)
  );
  not_cell not210 (
    .in (net262),
    .out (net271)
  );
  not_cell not211 (
    .in (net271),
    .out (net272)
  );
  not_cell not212 (
    .in (net272),
    .out (net273)
  );
  not_cell not213 (
    .in (net273),
    .out (net266)
  );
  not_cell not214 (
    .in (net274),
    .out (net275)
  );
  not_cell not215 (
    .in (net275),
    .out (net276)
  );
  not_cell not216 (
    .in (net276),
    .out (net277)
  );
  not_cell not217 (
    .in (net277),
    .out (net278)
  );
  not_cell not218 (
    .in (net270),
    .out (net279)
  );
  not_cell not219 (
    .in (net279),
    .out (net280)
  );
  not_cell not220 (
    .in (net280),
    .out (net281)
  );
  not_cell not221 (
    .in (net281),
    .out (net274)
  );
  not_cell not222 (
    .in (net282),
    .out (net283)
  );
  not_cell not223 (
    .in (net283),
    .out (net284)
  );
  not_cell not224 (
    .in (net284),
    .out (net285)
  );
  not_cell not225 (
    .in (net285),
    .out (net230)
  );
  not_cell not226 (
    .in (net278),
    .out (net286)
  );
  not_cell not227 (
    .in (net286),
    .out (net287)
  );
  not_cell not228 (
    .in (net287),
    .out (net288)
  );
  not_cell not229 (
    .in (net288),
    .out (net282)
  );
  not_cell not230 (
    .in (net289),
    .out (net290)
  );
  not_cell not231 (
    .in (net290),
    .out (net291)
  );
  not_cell not232 (
    .in (net291),
    .out (net292)
  );
  not_cell not233 (
    .in (net292),
    .out (net293)
  );
  not_cell not234 (
    .in (net294),
    .out (net295)
  );
  not_cell not235 (
    .in (net295),
    .out (net296)
  );
  not_cell not236 (
    .in (net296),
    .out (net297)
  );
  not_cell not237 (
    .in (net297),
    .out (net289)
  );
  not_cell not238 (
    .in (net298),
    .out (net299)
  );
  not_cell not239 (
    .in (net299),
    .out (net300)
  );
  not_cell not240 (
    .in (net300),
    .out (net301)
  );
  not_cell not241 (
    .in (net301),
    .out (net302)
  );
  not_cell not242 (
    .in (net293),
    .out (net303)
  );
  not_cell not243 (
    .in (net303),
    .out (net304)
  );
  not_cell not244 (
    .in (net304),
    .out (net305)
  );
  not_cell not245 (
    .in (net305),
    .out (net298)
  );
  not_cell not246 (
    .in (net306),
    .out (net307)
  );
  not_cell not247 (
    .in (net307),
    .out (net308)
  );
  not_cell not248 (
    .in (net308),
    .out (net309)
  );
  not_cell not249 (
    .in (net309),
    .out (net310)
  );
  not_cell not250 (
    .in (net302),
    .out (net311)
  );
  not_cell not251 (
    .in (net311),
    .out (net312)
  );
  not_cell not252 (
    .in (net312),
    .out (net313)
  );
  not_cell not253 (
    .in (net313),
    .out (net306)
  );
  not_cell not254 (
    .in (net314),
    .out (net315)
  );
  not_cell not255 (
    .in (net315),
    .out (net316)
  );
  not_cell not256 (
    .in (net316),
    .out (net317)
  );
  not_cell not257 (
    .in (net317),
    .out (net318)
  );
  not_cell not258 (
    .in (net310),
    .out (net319)
  );
  not_cell not259 (
    .in (net319),
    .out (net320)
  );
  not_cell not260 (
    .in (net320),
    .out (net321)
  );
  not_cell not261 (
    .in (net321),
    .out (net314)
  );
  not_cell not262 (
    .in (net322),
    .out (net323)
  );
  not_cell not263 (
    .in (net323),
    .out (net324)
  );
  not_cell not264 (
    .in (net324),
    .out (net325)
  );
  not_cell not265 (
    .in (net325),
    .out (net326)
  );
  not_cell not266 (
    .in (net254),
    .out (net327)
  );
  not_cell not267 (
    .in (net327),
    .out (net328)
  );
  not_cell not268 (
    .in (net328),
    .out (net329)
  );
  not_cell not269 (
    .in (net329),
    .out (net322)
  );
  not_cell not270 (
    .in (net330),
    .out (net331)
  );
  not_cell not271 (
    .in (net331),
    .out (net332)
  );
  not_cell not272 (
    .in (net332),
    .out (net333)
  );
  not_cell not273 (
    .in (net333),
    .out (net334)
  );
  not_cell not274 (
    .in (net326),
    .out (net335)
  );
  not_cell not275 (
    .in (net335),
    .out (net336)
  );
  not_cell not276 (
    .in (net336),
    .out (net337)
  );
  not_cell not277 (
    .in (net337),
    .out (net330)
  );
  not_cell not278 (
    .in (net338),
    .out (net339)
  );
  not_cell not279 (
    .in (net339),
    .out (net340)
  );
  not_cell not280 (
    .in (net340),
    .out (net341)
  );
  not_cell not281 (
    .in (net341),
    .out (net342)
  );
  not_cell not282 (
    .in (net334),
    .out (net343)
  );
  not_cell not283 (
    .in (net343),
    .out (net344)
  );
  not_cell not284 (
    .in (net344),
    .out (net345)
  );
  not_cell not285 (
    .in (net345),
    .out (net338)
  );
  not_cell not286 (
    .in (net346),
    .out (net347)
  );
  not_cell not287 (
    .in (net347),
    .out (net348)
  );
  not_cell not288 (
    .in (net348),
    .out (net349)
  );
  not_cell not289 (
    .in (net349),
    .out (net294)
  );
  not_cell not290 (
    .in (net342),
    .out (net350)
  );
  not_cell not291 (
    .in (net350),
    .out (net351)
  );
  not_cell not292 (
    .in (net351),
    .out (net352)
  );
  not_cell not293 (
    .in (net352),
    .out (net346)
  );
  not_cell not294 (
    .in (net353),
    .out (net354)
  );
  not_cell not295 (
    .in (net354),
    .out (net355)
  );
  not_cell not296 (
    .in (net355),
    .out (net356)
  );
  not_cell not297 (
    .in (net356),
    .out (net357)
  );
  not_cell not298 (
    .in (net358),
    .out (net359)
  );
  not_cell not299 (
    .in (net359),
    .out (net360)
  );
  not_cell not300 (
    .in (net360),
    .out (net361)
  );
  not_cell not301 (
    .in (net361),
    .out (net353)
  );
  not_cell not302 (
    .in (net362),
    .out (net363)
  );
  not_cell not303 (
    .in (net363),
    .out (net364)
  );
  not_cell not304 (
    .in (net364),
    .out (net365)
  );
  not_cell not305 (
    .in (net365),
    .out (net366)
  );
  not_cell not306 (
    .in (net357),
    .out (net367)
  );
  not_cell not307 (
    .in (net367),
    .out (net368)
  );
  not_cell not308 (
    .in (net368),
    .out (net369)
  );
  not_cell not309 (
    .in (net369),
    .out (net362)
  );
  not_cell not310 (
    .in (net370),
    .out (net371)
  );
  not_cell not311 (
    .in (net371),
    .out (net372)
  );
  not_cell not312 (
    .in (net372),
    .out (net373)
  );
  not_cell not313 (
    .in (net373),
    .out (net374)
  );
  not_cell not314 (
    .in (net366),
    .out (net375)
  );
  not_cell not315 (
    .in (net375),
    .out (net376)
  );
  not_cell not316 (
    .in (net376),
    .out (net377)
  );
  not_cell not317 (
    .in (net377),
    .out (net370)
  );
  not_cell not318 (
    .in (net378),
    .out (net379)
  );
  not_cell not319 (
    .in (net379),
    .out (net380)
  );
  not_cell not320 (
    .in (net380),
    .out (net381)
  );
  not_cell not321 (
    .in (net381),
    .out (net382)
  );
  not_cell not322 (
    .in (net374),
    .out (net383)
  );
  not_cell not323 (
    .in (net383),
    .out (net384)
  );
  not_cell not324 (
    .in (net384),
    .out (net385)
  );
  not_cell not325 (
    .in (net385),
    .out (net378)
  );
  not_cell not326 (
    .in (net386),
    .out (net387)
  );
  not_cell not327 (
    .in (net387),
    .out (net388)
  );
  not_cell not328 (
    .in (net388),
    .out (net389)
  );
  not_cell not329 (
    .in (net389),
    .out (net390)
  );
  not_cell not330 (
    .in (net318),
    .out (net391)
  );
  not_cell not331 (
    .in (net391),
    .out (net392)
  );
  not_cell not332 (
    .in (net392),
    .out (net393)
  );
  not_cell not333 (
    .in (net393),
    .out (net386)
  );
  not_cell not334 (
    .in (net394),
    .out (net395)
  );
  not_cell not335 (
    .in (net395),
    .out (net396)
  );
  not_cell not336 (
    .in (net396),
    .out (net397)
  );
  not_cell not337 (
    .in (net397),
    .out (net398)
  );
  not_cell not338 (
    .in (net390),
    .out (net399)
  );
  not_cell not339 (
    .in (net399),
    .out (net400)
  );
  not_cell not340 (
    .in (net400),
    .out (net401)
  );
  not_cell not341 (
    .in (net401),
    .out (net394)
  );
  not_cell not342 (
    .in (net402),
    .out (net403)
  );
  not_cell not343 (
    .in (net403),
    .out (net404)
  );
  not_cell not344 (
    .in (net404),
    .out (net405)
  );
  not_cell not345 (
    .in (net405),
    .out (net406)
  );
  not_cell not346 (
    .in (net398),
    .out (net407)
  );
  not_cell not347 (
    .in (net407),
    .out (net408)
  );
  not_cell not348 (
    .in (net408),
    .out (net409)
  );
  not_cell not349 (
    .in (net409),
    .out (net402)
  );
  not_cell not350 (
    .in (net410),
    .out (net411)
  );
  not_cell not351 (
    .in (net411),
    .out (net412)
  );
  not_cell not352 (
    .in (net412),
    .out (net413)
  );
  not_cell not353 (
    .in (net413),
    .out (net358)
  );
  not_cell not354 (
    .in (net406),
    .out (net414)
  );
  not_cell not355 (
    .in (net414),
    .out (net415)
  );
  not_cell not356 (
    .in (net415),
    .out (net416)
  );
  not_cell not357 (
    .in (net416),
    .out (net410)
  );
  not_cell not358 (
    .in (net417),
    .out (net418)
  );
  not_cell not359 (
    .in (net418),
    .out (net419)
  );
  not_cell not360 (
    .in (net419),
    .out (net420)
  );
  not_cell not361 (
    .in (net420),
    .out (net421)
  );
  not_cell not362 (
    .in (net422),
    .out (net423)
  );
  not_cell not363 (
    .in (net423),
    .out (net424)
  );
  not_cell not364 (
    .in (net424),
    .out (net425)
  );
  not_cell not365 (
    .in (net425),
    .out (net417)
  );
  not_cell not366 (
    .in (net426),
    .out (net427)
  );
  not_cell not367 (
    .in (net427),
    .out (net428)
  );
  not_cell not368 (
    .in (net428),
    .out (net429)
  );
  not_cell not369 (
    .in (net429),
    .out (net430)
  );
  not_cell not370 (
    .in (net421),
    .out (net431)
  );
  not_cell not371 (
    .in (net431),
    .out (net432)
  );
  not_cell not372 (
    .in (net432),
    .out (net433)
  );
  not_cell not373 (
    .in (net433),
    .out (net426)
  );
  not_cell not374 (
    .in (net434),
    .out (net435)
  );
  not_cell not375 (
    .in (net435),
    .out (net436)
  );
  not_cell not376 (
    .in (net436),
    .out (net437)
  );
  not_cell not377 (
    .in (net437),
    .out (net438)
  );
  not_cell not378 (
    .in (net430),
    .out (net439)
  );
  not_cell not379 (
    .in (net439),
    .out (net440)
  );
  not_cell not380 (
    .in (net440),
    .out (net441)
  );
  not_cell not381 (
    .in (net441),
    .out (net434)
  );
  not_cell not382 (
    .in (net442),
    .out (net443)
  );
  not_cell not383 (
    .in (net443),
    .out (net444)
  );
  not_cell not384 (
    .in (net444),
    .out (net445)
  );
  not_cell not385 (
    .in (net445),
    .out (net446)
  );
  not_cell not386 (
    .in (net438),
    .out (net447)
  );
  not_cell not387 (
    .in (net447),
    .out (net448)
  );
  not_cell not388 (
    .in (net448),
    .out (net449)
  );
  not_cell not389 (
    .in (net449),
    .out (net442)
  );
  not_cell not390 (
    .in (net450),
    .out (net451)
  );
  not_cell not391 (
    .in (net451),
    .out (net452)
  );
  not_cell not392 (
    .in (net452),
    .out (net453)
  );
  not_cell not393 (
    .in (net453),
    .out (net454)
  );
  not_cell not394 (
    .in (net382),
    .out (net455)
  );
  not_cell not395 (
    .in (net455),
    .out (net456)
  );
  not_cell not396 (
    .in (net456),
    .out (net457)
  );
  not_cell not397 (
    .in (net457),
    .out (net450)
  );
  not_cell not398 (
    .in (net458),
    .out (net459)
  );
  not_cell not399 (
    .in (net459),
    .out (net460)
  );
  not_cell not400 (
    .in (net460),
    .out (net461)
  );
  not_cell not401 (
    .in (net461),
    .out (net462)
  );
  not_cell not402 (
    .in (net454),
    .out (net463)
  );
  not_cell not403 (
    .in (net463),
    .out (net464)
  );
  not_cell not404 (
    .in (net464),
    .out (net465)
  );
  not_cell not405 (
    .in (net465),
    .out (net458)
  );
  not_cell not406 (
    .in (net466),
    .out (net467)
  );
  not_cell not407 (
    .in (net467),
    .out (net468)
  );
  not_cell not408 (
    .in (net468),
    .out (net469)
  );
  not_cell not409 (
    .in (net469),
    .out (net470)
  );
  not_cell not410 (
    .in (net462),
    .out (net471)
  );
  not_cell not411 (
    .in (net471),
    .out (net472)
  );
  not_cell not412 (
    .in (net472),
    .out (net473)
  );
  not_cell not413 (
    .in (net473),
    .out (net466)
  );
  not_cell not414 (
    .in (net474),
    .out (net475)
  );
  not_cell not415 (
    .in (net475),
    .out (net476)
  );
  not_cell not416 (
    .in (net476),
    .out (net477)
  );
  not_cell not417 (
    .in (net477),
    .out (net422)
  );
  not_cell not418 (
    .in (net470),
    .out (net478)
  );
  not_cell not419 (
    .in (net478),
    .out (net479)
  );
  not_cell not420 (
    .in (net479),
    .out (net480)
  );
  not_cell not421 (
    .in (net480),
    .out (net474)
  );
  or_cell or1 (
    .a (net11),
    .b (net446),
    .out (net4)
  );
endmodule
