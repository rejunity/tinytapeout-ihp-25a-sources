(* blackbox *) (* keep *)
module my_logo ();
endmodule
