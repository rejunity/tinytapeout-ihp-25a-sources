/* Automatically generated from https://wokwi.com/projects/413921288682183681 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_413921288682183681(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = ui_in[0];
  wire net3 = ui_in[1];
  wire net4 = ui_in[2];
  wire net5 = ui_in[3];
  wire net6 = ui_in[4];
  wire net7 = ui_in[5];
  wire net8 = ui_in[6];
  wire net9 = ui_in[7];
  wire net10;
  wire net11;
  wire net12;
  wire net13 = 1'b1;
  wire net14 = 1'b1;
  wire net15 = 1'b0;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26 = 1'b0;

  assign uo_out[0] = net10;
  assign uo_out[1] = net11;
  assign uo_out[2] = net12;
  assign uo_out[3] = net9;
  assign uo_out[4] = net1;
  assign uo_out[5] = 0;
  assign uo_out[6] = 0;
  assign uo_out[7] = 0;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  or_cell or1 (
    .a (net2),
    .b (net4),
    .out (net17)
  );
  or_cell or2 (
    .a (net6),
    .b (net8),
    .out (net18)
  );
  or_cell or3 (
    .a (net3),
    .b (net4),
    .out (net19)
  );
  or_cell or4 (
    .a (net7),
    .b (net8),
    .out (net20)
  );
  or_cell or5 (
    .a (net5),
    .b (net6),
    .out (net21)
  );
  or_cell or6 (
    .a (net7),
    .b (net8),
    .out (net22)
  );
  or_cell or7 (
    .a (net17),
    .b (net18),
    .out (net23)
  );
  or_cell or8 (
    .a (net19),
    .b (net20),
    .out (net24)
  );
  or_cell or9 (
    .a (net21),
    .b (net22),
    .out (net25)
  );
  xor_cell xor1 (
    .a (net23),
    .b (net9),
    .out (net10)
  );
  xor_cell xor2 (
    .a (net24),
    .b (net9),
    .out (net11)
  );
  xor_cell xor3 (
    .a (net25),
    .b (net9),
    .out (net12)
  );
endmodule
