VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 109.900 BY 20.300 ;
  OBS
      LAYER met1 ;
        RECT 0.000 19.950 8.050 20.300 ;
      LAYER met1 ;
        RECT 8.050 19.950 11.550 20.300 ;
      LAYER met1 ;
        RECT 11.550 19.950 22.050 20.300 ;
      LAYER met1 ;
        RECT 22.050 19.950 24.500 20.300 ;
      LAYER met1 ;
        RECT 24.500 19.950 31.500 20.300 ;
      LAYER met1 ;
        RECT 31.500 19.950 33.950 20.300 ;
      LAYER met1 ;
        RECT 33.950 19.950 54.250 20.300 ;
      LAYER met1 ;
        RECT 54.250 19.950 56.700 20.300 ;
      LAYER met1 ;
        RECT 56.700 19.950 68.950 20.300 ;
      LAYER met1 ;
        RECT 68.950 19.950 71.050 20.300 ;
      LAYER met1 ;
        RECT 71.050 19.950 109.900 20.300 ;
        RECT 0.000 19.600 6.650 19.950 ;
      LAYER met1 ;
        RECT 6.650 19.600 12.950 19.950 ;
      LAYER met1 ;
        RECT 12.950 19.600 21.700 19.950 ;
      LAYER met1 ;
        RECT 21.700 19.600 24.500 19.950 ;
      LAYER met1 ;
        RECT 24.500 19.600 30.450 19.950 ;
      LAYER met1 ;
        RECT 30.450 19.600 35.000 19.950 ;
      LAYER met1 ;
        RECT 35.000 19.600 42.700 19.950 ;
      LAYER met1 ;
        RECT 42.700 19.600 45.500 19.950 ;
      LAYER met1 ;
        RECT 45.500 19.600 48.650 19.950 ;
      LAYER met1 ;
        RECT 48.650 19.600 51.100 19.950 ;
      LAYER met1 ;
        RECT 51.100 19.600 53.550 19.950 ;
      LAYER met1 ;
        RECT 53.550 19.600 57.400 19.950 ;
      LAYER met1 ;
        RECT 57.400 19.600 58.800 19.950 ;
      LAYER met1 ;
        RECT 58.800 19.600 61.950 19.950 ;
      LAYER met1 ;
        RECT 61.950 19.600 67.900 19.950 ;
      LAYER met1 ;
        RECT 67.900 19.600 72.100 19.950 ;
      LAYER met1 ;
        RECT 72.100 19.600 86.450 19.950 ;
      LAYER met1 ;
        RECT 86.450 19.600 92.050 19.950 ;
      LAYER met1 ;
        RECT 92.050 19.600 109.900 19.950 ;
        RECT 0.000 19.250 5.600 19.600 ;
      LAYER met1 ;
        RECT 5.600 19.250 13.650 19.600 ;
      LAYER met1 ;
        RECT 13.650 19.250 21.000 19.600 ;
      LAYER met1 ;
        RECT 21.000 19.250 24.500 19.600 ;
      LAYER met1 ;
        RECT 24.500 19.250 30.100 19.600 ;
      LAYER met1 ;
        RECT 30.100 19.250 32.200 19.600 ;
      LAYER met1 ;
        RECT 32.200 19.250 33.250 19.600 ;
      LAYER met1 ;
        RECT 33.250 19.250 35.350 19.600 ;
      LAYER met1 ;
        RECT 35.350 19.250 43.400 19.600 ;
        RECT 0.000 18.900 4.900 19.250 ;
      LAYER met1 ;
        RECT 4.900 18.900 14.350 19.250 ;
      LAYER met1 ;
        RECT 14.350 18.900 20.300 19.250 ;
      LAYER met1 ;
        RECT 20.300 18.900 24.500 19.250 ;
      LAYER met1 ;
        RECT 24.500 18.900 29.750 19.250 ;
      LAYER met1 ;
        RECT 29.750 18.900 31.850 19.250 ;
      LAYER met1 ;
        RECT 31.850 18.900 33.600 19.250 ;
      LAYER met1 ;
        RECT 33.600 18.900 35.700 19.250 ;
      LAYER met1 ;
        RECT 35.700 18.900 43.400 19.250 ;
      LAYER met1 ;
        RECT 43.400 18.900 44.800 19.600 ;
      LAYER met1 ;
        RECT 44.800 18.900 49.350 19.600 ;
      LAYER met1 ;
        RECT 49.350 19.250 50.400 19.600 ;
      LAYER met1 ;
        RECT 50.400 19.250 53.200 19.600 ;
      LAYER met1 ;
        RECT 53.200 19.250 54.250 19.600 ;
      LAYER met1 ;
        RECT 54.250 19.250 55.650 19.600 ;
      LAYER met1 ;
        RECT 55.650 19.250 57.400 19.600 ;
      LAYER met1 ;
        RECT 57.400 19.250 59.500 19.600 ;
      LAYER met1 ;
        RECT 59.500 19.250 61.250 19.600 ;
      LAYER met1 ;
        RECT 61.250 19.250 67.550 19.600 ;
      LAYER met1 ;
        RECT 67.550 19.250 68.950 19.600 ;
      LAYER met1 ;
        RECT 68.950 19.250 70.000 19.600 ;
      LAYER met1 ;
        RECT 70.000 19.250 72.100 19.600 ;
      LAYER met1 ;
        RECT 0.000 18.550 4.550 18.900 ;
      LAYER met1 ;
        RECT 4.550 18.550 8.750 18.900 ;
      LAYER met1 ;
        RECT 8.750 18.550 10.850 18.900 ;
      LAYER met1 ;
        RECT 10.850 18.550 15.050 18.900 ;
      LAYER met1 ;
        RECT 15.050 18.550 19.950 18.900 ;
      LAYER met1 ;
        RECT 19.950 18.550 21.700 18.900 ;
      LAYER met1 ;
        RECT 21.700 18.550 22.050 18.900 ;
        RECT 0.000 18.200 3.850 18.550 ;
      LAYER met1 ;
        RECT 3.850 18.200 7.000 18.550 ;
      LAYER met1 ;
        RECT 7.000 18.200 12.250 18.550 ;
      LAYER met1 ;
        RECT 12.250 18.200 15.400 18.550 ;
      LAYER met1 ;
        RECT 15.400 18.200 19.950 18.550 ;
      LAYER met1 ;
        RECT 19.950 18.200 21.000 18.550 ;
      LAYER met1 ;
        RECT 21.000 18.200 22.050 18.550 ;
        RECT 0.000 17.850 3.500 18.200 ;
      LAYER met1 ;
        RECT 3.500 17.850 6.300 18.200 ;
      LAYER met1 ;
        RECT 6.300 17.850 13.300 18.200 ;
      LAYER met1 ;
        RECT 13.300 17.850 16.100 18.200 ;
      LAYER met1 ;
        RECT 16.100 17.850 19.950 18.200 ;
      LAYER met1 ;
        RECT 19.950 17.850 20.300 18.200 ;
      LAYER met1 ;
        RECT 20.300 17.850 22.050 18.200 ;
        RECT 0.000 17.500 3.150 17.850 ;
      LAYER met1 ;
        RECT 3.150 17.500 5.600 17.850 ;
      LAYER met1 ;
        RECT 5.600 17.500 14.000 17.850 ;
      LAYER met1 ;
        RECT 14.000 17.500 16.450 17.850 ;
      LAYER met1 ;
        RECT 16.450 17.500 22.050 17.850 ;
        RECT 0.000 17.150 2.800 17.500 ;
      LAYER met1 ;
        RECT 2.800 17.150 4.900 17.500 ;
      LAYER met1 ;
        RECT 4.900 17.150 14.350 17.500 ;
      LAYER met1 ;
        RECT 14.350 17.150 16.800 17.500 ;
      LAYER met1 ;
        RECT 16.800 17.150 22.050 17.500 ;
        RECT 0.000 16.800 2.450 17.150 ;
      LAYER met1 ;
        RECT 2.450 16.800 4.550 17.150 ;
      LAYER met1 ;
        RECT 4.550 16.800 15.050 17.150 ;
      LAYER met1 ;
        RECT 15.050 16.800 17.150 17.150 ;
      LAYER met1 ;
        RECT 17.150 16.800 22.050 17.150 ;
        RECT 0.000 16.450 2.100 16.800 ;
      LAYER met1 ;
        RECT 2.100 16.450 4.200 16.800 ;
      LAYER met1 ;
        RECT 4.200 16.450 15.400 16.800 ;
      LAYER met1 ;
        RECT 15.400 16.450 17.500 16.800 ;
      LAYER met1 ;
        RECT 0.000 15.750 1.750 16.450 ;
      LAYER met1 ;
        RECT 1.750 16.100 3.850 16.450 ;
      LAYER met1 ;
        RECT 3.850 16.100 15.750 16.450 ;
      LAYER met1 ;
        RECT 15.750 16.100 17.500 16.450 ;
      LAYER met1 ;
        RECT 17.500 16.100 22.050 16.800 ;
      LAYER met1 ;
        RECT 1.750 15.750 11.550 16.100 ;
      LAYER met1 ;
        RECT 11.550 15.750 16.100 16.100 ;
      LAYER met1 ;
        RECT 16.100 15.750 17.850 16.100 ;
      LAYER met1 ;
        RECT 17.850 15.750 22.050 16.100 ;
        RECT 0.000 15.050 1.400 15.750 ;
      LAYER met1 ;
        RECT 1.400 15.050 11.550 15.750 ;
      LAYER met1 ;
        RECT 11.550 15.050 16.450 15.750 ;
      LAYER met1 ;
        RECT 16.450 15.050 18.200 15.750 ;
      LAYER met1 ;
        RECT 18.200 15.050 22.050 15.750 ;
        RECT 0.000 14.350 1.050 15.050 ;
      LAYER met1 ;
        RECT 1.050 14.350 11.550 15.050 ;
      LAYER met1 ;
        RECT 11.550 14.350 16.800 15.050 ;
      LAYER met1 ;
        RECT 16.800 14.350 18.550 15.050 ;
      LAYER met1 ;
        RECT 18.550 14.350 22.050 15.050 ;
        RECT 0.000 13.650 0.700 14.350 ;
      LAYER met1 ;
        RECT 0.700 13.650 11.550 14.350 ;
      LAYER met1 ;
        RECT 11.550 13.650 17.150 14.350 ;
      LAYER met1 ;
        RECT 17.150 13.650 18.900 14.350 ;
      LAYER met1 ;
        RECT 0.000 13.300 5.600 13.650 ;
      LAYER met1 ;
        RECT 5.600 13.300 8.750 13.650 ;
      LAYER met1 ;
        RECT 0.000 12.600 5.950 13.300 ;
        RECT 0.000 12.250 0.350 12.600 ;
      LAYER met1 ;
        RECT 0.350 12.250 1.750 12.600 ;
        RECT 0.000 11.550 1.750 12.250 ;
      LAYER met1 ;
        RECT 1.750 11.550 5.950 12.600 ;
      LAYER met1 ;
        RECT 0.000 9.450 1.400 11.550 ;
      LAYER met1 ;
        RECT 1.400 9.450 5.950 11.550 ;
      LAYER met1 ;
        RECT 5.950 11.200 8.750 13.300 ;
      LAYER met1 ;
        RECT 8.750 12.950 17.500 13.650 ;
      LAYER met1 ;
        RECT 17.500 13.300 18.900 13.650 ;
      LAYER met1 ;
        RECT 18.900 13.300 22.050 14.350 ;
      LAYER met1 ;
        RECT 17.500 12.950 19.250 13.300 ;
      LAYER met1 ;
        RECT 8.750 11.200 17.850 12.950 ;
      LAYER met1 ;
        RECT 17.850 11.900 19.250 12.950 ;
      LAYER met1 ;
        RECT 19.250 11.900 22.050 13.300 ;
      LAYER met1 ;
        RECT 0.000 8.750 1.750 9.450 ;
      LAYER met1 ;
        RECT 0.000 7.350 0.350 8.750 ;
      LAYER met1 ;
        RECT 0.350 7.700 1.750 8.750 ;
      LAYER met1 ;
        RECT 1.750 7.700 5.950 9.450 ;
      LAYER met1 ;
        RECT 5.950 8.750 16.100 11.200 ;
      LAYER met1 ;
        RECT 16.100 8.750 17.850 11.200 ;
      LAYER met1 ;
        RECT 17.850 9.100 19.600 11.900 ;
      LAYER met1 ;
        RECT 19.600 10.850 22.050 11.900 ;
      LAYER met1 ;
        RECT 22.050 10.850 24.500 18.900 ;
      LAYER met1 ;
        RECT 24.500 18.200 29.400 18.900 ;
      LAYER met1 ;
        RECT 29.400 18.200 31.500 18.900 ;
      LAYER met1 ;
        RECT 24.500 17.500 29.050 18.200 ;
      LAYER met1 ;
        RECT 29.050 17.500 31.500 18.200 ;
      LAYER met1 ;
        RECT 24.500 12.600 28.700 17.500 ;
      LAYER met1 ;
        RECT 28.700 16.450 31.500 17.500 ;
      LAYER met1 ;
        RECT 31.500 16.450 33.950 18.900 ;
      LAYER met1 ;
        RECT 33.950 18.200 36.050 18.900 ;
      LAYER met1 ;
        RECT 36.050 18.200 43.750 18.900 ;
      LAYER met1 ;
        RECT 43.750 18.200 45.150 18.900 ;
      LAYER met1 ;
        RECT 45.150 18.550 49.350 18.900 ;
      LAYER met1 ;
        RECT 49.350 18.550 50.050 19.250 ;
      LAYER met1 ;
        RECT 50.050 18.900 52.850 19.250 ;
      LAYER met1 ;
        RECT 52.850 18.900 53.900 19.250 ;
      LAYER met1 ;
        RECT 53.900 18.900 56.000 19.250 ;
      LAYER met1 ;
        RECT 56.000 18.900 57.400 19.250 ;
      LAYER met1 ;
        RECT 57.400 18.900 59.850 19.250 ;
      LAYER met1 ;
        RECT 33.950 17.500 36.400 18.200 ;
      LAYER met1 ;
        RECT 36.400 17.500 44.100 18.200 ;
      LAYER met1 ;
        RECT 44.100 17.850 45.150 18.200 ;
      LAYER met1 ;
        RECT 45.150 17.850 49.000 18.550 ;
      LAYER met1 ;
        RECT 49.000 18.200 50.050 18.550 ;
      LAYER met1 ;
        RECT 50.050 18.200 52.500 18.900 ;
      LAYER met1 ;
        RECT 49.000 17.850 49.700 18.200 ;
        RECT 28.700 13.650 31.150 16.450 ;
      LAYER met1 ;
        RECT 31.150 13.650 33.950 16.450 ;
      LAYER met1 ;
        RECT 28.700 12.600 31.500 13.650 ;
      LAYER met1 ;
        RECT 24.500 11.550 29.050 12.600 ;
      LAYER met1 ;
        RECT 29.050 11.550 31.500 12.600 ;
      LAYER met1 ;
        RECT 24.500 11.200 29.400 11.550 ;
      LAYER met1 ;
        RECT 29.400 11.200 31.500 11.550 ;
      LAYER met1 ;
        RECT 31.500 11.200 33.950 13.650 ;
      LAYER met1 ;
        RECT 33.950 12.600 36.750 17.500 ;
      LAYER met1 ;
        RECT 36.750 17.150 44.100 17.500 ;
      LAYER met1 ;
        RECT 44.100 17.150 45.500 17.850 ;
      LAYER met1 ;
        RECT 36.750 16.100 44.450 17.150 ;
      LAYER met1 ;
        RECT 44.450 16.800 45.500 17.150 ;
      LAYER met1 ;
        RECT 45.500 16.800 48.650 17.850 ;
      LAYER met1 ;
        RECT 48.650 17.150 49.700 17.850 ;
      LAYER met1 ;
        RECT 49.700 17.150 52.500 18.200 ;
      LAYER met1 ;
        RECT 52.500 17.850 53.550 18.900 ;
      LAYER met1 ;
        RECT 53.550 18.550 56.350 18.900 ;
      LAYER met1 ;
        RECT 56.350 18.550 57.050 18.900 ;
      LAYER met1 ;
        RECT 57.050 18.550 59.850 18.900 ;
        RECT 53.550 17.850 59.850 18.550 ;
      LAYER met1 ;
        RECT 52.500 17.500 53.900 17.850 ;
      LAYER met1 ;
        RECT 53.900 17.500 59.850 17.850 ;
      LAYER met1 ;
        RECT 52.500 17.150 54.250 17.500 ;
      LAYER met1 ;
        RECT 54.250 17.150 59.850 17.500 ;
      LAYER met1 ;
        RECT 48.650 16.800 49.350 17.150 ;
      LAYER met1 ;
        RECT 49.350 16.800 52.850 17.150 ;
      LAYER met1 ;
        RECT 52.850 16.800 54.950 17.150 ;
      LAYER met1 ;
        RECT 54.950 16.800 59.850 17.150 ;
      LAYER met1 ;
        RECT 44.450 16.100 45.850 16.800 ;
      LAYER met1 ;
        RECT 45.850 16.100 48.300 16.800 ;
      LAYER met1 ;
        RECT 48.300 16.100 49.350 16.800 ;
      LAYER met1 ;
        RECT 49.350 16.450 53.200 16.800 ;
      LAYER met1 ;
        RECT 53.200 16.450 55.650 16.800 ;
      LAYER met1 ;
        RECT 55.650 16.450 59.850 16.800 ;
        RECT 49.350 16.100 53.550 16.450 ;
      LAYER met1 ;
        RECT 53.550 16.100 56.350 16.450 ;
      LAYER met1 ;
        RECT 56.350 16.100 59.850 16.450 ;
        RECT 36.750 15.400 44.800 16.100 ;
      LAYER met1 ;
        RECT 44.800 15.400 46.200 16.100 ;
      LAYER met1 ;
        RECT 46.200 15.750 48.300 16.100 ;
      LAYER met1 ;
        RECT 48.300 15.750 49.000 16.100 ;
      LAYER met1 ;
        RECT 49.000 15.750 53.900 16.100 ;
      LAYER met1 ;
        RECT 53.900 15.750 56.700 16.100 ;
      LAYER met1 ;
        RECT 56.700 15.750 59.850 16.100 ;
        RECT 36.750 14.350 45.150 15.400 ;
      LAYER met1 ;
        RECT 45.150 15.050 46.200 15.400 ;
      LAYER met1 ;
        RECT 46.200 15.050 47.950 15.750 ;
      LAYER met1 ;
        RECT 47.950 15.050 49.000 15.750 ;
      LAYER met1 ;
        RECT 49.000 15.400 54.600 15.750 ;
      LAYER met1 ;
        RECT 54.600 15.400 57.050 15.750 ;
      LAYER met1 ;
        RECT 57.050 15.400 59.850 15.750 ;
        RECT 49.000 15.050 55.300 15.400 ;
      LAYER met1 ;
        RECT 55.300 15.050 57.400 15.400 ;
      LAYER met1 ;
        RECT 57.400 15.050 59.850 15.400 ;
      LAYER met1 ;
        RECT 45.150 14.350 46.550 15.050 ;
      LAYER met1 ;
        RECT 46.550 14.700 47.950 15.050 ;
      LAYER met1 ;
        RECT 47.950 14.700 48.650 15.050 ;
      LAYER met1 ;
        RECT 48.650 14.700 56.000 15.050 ;
      LAYER met1 ;
        RECT 56.000 14.700 57.750 15.050 ;
      LAYER met1 ;
        RECT 36.750 13.300 45.500 14.350 ;
      LAYER met1 ;
        RECT 45.500 14.000 46.550 14.350 ;
      LAYER met1 ;
        RECT 46.550 14.000 47.600 14.700 ;
      LAYER met1 ;
        RECT 47.600 14.350 48.650 14.700 ;
      LAYER met1 ;
        RECT 48.650 14.350 56.350 14.700 ;
      LAYER met1 ;
        RECT 56.350 14.350 57.750 14.700 ;
        RECT 45.500 13.300 46.900 14.000 ;
      LAYER met1 ;
        RECT 46.900 13.650 47.600 14.000 ;
      LAYER met1 ;
        RECT 47.600 13.650 48.300 14.350 ;
      LAYER met1 ;
        RECT 48.300 13.650 56.700 14.350 ;
        RECT 46.900 13.300 47.250 13.650 ;
      LAYER met1 ;
        RECT 47.250 13.300 48.300 13.650 ;
      LAYER met1 ;
        RECT 48.300 13.300 52.500 13.650 ;
      LAYER met1 ;
        RECT 52.500 13.300 52.850 13.650 ;
      LAYER met1 ;
        RECT 52.850 13.300 56.700 13.650 ;
        RECT 36.750 12.600 45.850 13.300 ;
      LAYER met1 ;
        RECT 45.850 12.600 47.950 13.300 ;
        RECT 33.950 11.900 36.400 12.600 ;
      LAYER met1 ;
        RECT 36.400 11.900 46.200 12.600 ;
      LAYER met1 ;
        RECT 46.200 12.250 47.950 12.600 ;
      LAYER met1 ;
        RECT 47.950 12.250 52.500 13.300 ;
      LAYER met1 ;
        RECT 52.500 12.950 53.200 13.300 ;
      LAYER met1 ;
        RECT 53.200 12.950 56.700 13.300 ;
      LAYER met1 ;
        RECT 56.700 12.950 57.750 14.350 ;
      LAYER met1 ;
        RECT 57.750 12.950 59.850 15.050 ;
      LAYER met1 ;
        RECT 52.500 12.600 53.550 12.950 ;
      LAYER met1 ;
        RECT 53.550 12.600 56.350 12.950 ;
      LAYER met1 ;
        RECT 56.350 12.600 57.400 12.950 ;
        RECT 52.500 12.250 53.900 12.600 ;
      LAYER met1 ;
        RECT 53.900 12.250 56.000 12.600 ;
      LAYER met1 ;
        RECT 56.000 12.250 57.400 12.600 ;
      LAYER met1 ;
        RECT 57.400 12.250 59.850 12.950 ;
      LAYER met1 ;
        RECT 59.850 12.600 60.900 19.250 ;
      LAYER met1 ;
        RECT 60.900 18.900 67.200 19.250 ;
      LAYER met1 ;
        RECT 67.200 18.900 68.250 19.250 ;
      LAYER met1 ;
        RECT 68.250 18.900 70.700 19.250 ;
      LAYER met1 ;
        RECT 70.700 18.900 72.100 19.250 ;
      LAYER met1 ;
        RECT 72.100 18.900 79.100 19.600 ;
        RECT 60.900 18.550 66.850 18.900 ;
      LAYER met1 ;
        RECT 66.850 18.550 67.900 18.900 ;
      LAYER met1 ;
        RECT 67.900 18.550 71.400 18.900 ;
      LAYER met1 ;
        RECT 71.400 18.550 71.750 18.900 ;
      LAYER met1 ;
        RECT 71.750 18.550 79.100 18.900 ;
        RECT 60.900 17.850 66.500 18.550 ;
      LAYER met1 ;
        RECT 66.500 17.850 67.550 18.550 ;
      LAYER met1 ;
        RECT 67.550 18.200 79.100 18.550 ;
      LAYER met1 ;
        RECT 79.100 18.200 85.400 19.600 ;
      LAYER met1 ;
        RECT 85.400 18.200 86.100 19.600 ;
      LAYER met1 ;
        RECT 86.100 18.200 92.050 19.600 ;
      LAYER met1 ;
        RECT 92.050 18.200 93.100 19.600 ;
        RECT 67.550 17.850 83.300 18.200 ;
        RECT 60.900 17.150 66.150 17.850 ;
      LAYER met1 ;
        RECT 66.150 17.150 67.200 17.850 ;
      LAYER met1 ;
        RECT 60.900 14.000 65.800 17.150 ;
      LAYER met1 ;
        RECT 65.800 14.000 67.200 17.150 ;
      LAYER met1 ;
        RECT 67.200 14.000 83.300 17.850 ;
        RECT 60.900 13.300 66.150 14.000 ;
      LAYER met1 ;
        RECT 66.150 13.300 67.550 14.000 ;
      LAYER met1 ;
        RECT 67.550 13.650 83.300 14.000 ;
        RECT 67.550 13.300 79.100 13.650 ;
        RECT 60.900 12.950 64.750 13.300 ;
      LAYER met1 ;
        RECT 64.750 12.950 65.100 13.300 ;
      LAYER met1 ;
        RECT 65.100 12.950 66.150 13.300 ;
      LAYER met1 ;
        RECT 66.150 12.950 67.900 13.300 ;
      LAYER met1 ;
        RECT 67.900 12.950 79.100 13.300 ;
        RECT 60.900 12.600 64.400 12.950 ;
      LAYER met1 ;
        RECT 59.850 12.250 61.250 12.600 ;
      LAYER met1 ;
        RECT 61.250 12.250 64.400 12.600 ;
      LAYER met1 ;
        RECT 64.400 12.250 65.100 12.950 ;
      LAYER met1 ;
        RECT 65.100 12.600 66.500 12.950 ;
      LAYER met1 ;
        RECT 66.500 12.600 68.250 12.950 ;
      LAYER met1 ;
        RECT 68.250 12.600 71.400 12.950 ;
      LAYER met1 ;
        RECT 71.400 12.600 72.450 12.950 ;
      LAYER met1 ;
        RECT 72.450 12.600 79.100 12.950 ;
        RECT 65.100 12.250 66.850 12.600 ;
      LAYER met1 ;
        RECT 66.850 12.250 68.600 12.600 ;
      LAYER met1 ;
        RECT 68.600 12.250 71.050 12.600 ;
      LAYER met1 ;
        RECT 71.050 12.250 72.100 12.600 ;
      LAYER met1 ;
        RECT 72.100 12.250 79.100 12.600 ;
      LAYER met1 ;
        RECT 33.950 11.200 36.050 11.900 ;
      LAYER met1 ;
        RECT 36.050 11.550 46.200 11.900 ;
      LAYER met1 ;
        RECT 46.200 11.550 47.600 12.250 ;
      LAYER met1 ;
        RECT 47.600 11.900 52.500 12.250 ;
      LAYER met1 ;
        RECT 52.500 11.900 54.600 12.250 ;
      LAYER met1 ;
        RECT 54.600 11.900 55.300 12.250 ;
      LAYER met1 ;
        RECT 55.300 11.900 57.050 12.250 ;
      LAYER met1 ;
        RECT 57.050 11.900 59.500 12.250 ;
      LAYER met1 ;
        RECT 59.500 11.900 62.300 12.250 ;
      LAYER met1 ;
        RECT 62.300 11.900 63.350 12.250 ;
      LAYER met1 ;
        RECT 63.350 11.900 65.100 12.250 ;
      LAYER met1 ;
        RECT 65.100 11.900 67.200 12.250 ;
      LAYER met1 ;
        RECT 67.200 11.900 71.750 12.250 ;
      LAYER met1 ;
        RECT 71.750 11.900 79.100 12.250 ;
        RECT 47.600 11.550 52.850 11.900 ;
      LAYER met1 ;
        RECT 52.850 11.550 56.700 11.900 ;
      LAYER met1 ;
        RECT 56.700 11.550 58.800 11.900 ;
        RECT 36.050 11.200 46.550 11.550 ;
      LAYER met1 ;
        RECT 46.550 11.200 47.250 11.550 ;
      LAYER met1 ;
        RECT 47.250 11.200 53.550 11.550 ;
      LAYER met1 ;
        RECT 53.550 11.200 56.000 11.550 ;
      LAYER met1 ;
        RECT 56.000 11.200 58.800 11.550 ;
      LAYER met1 ;
        RECT 58.800 11.200 64.750 11.900 ;
      LAYER met1 ;
        RECT 64.750 11.550 67.550 11.900 ;
      LAYER met1 ;
        RECT 67.550 11.550 71.050 11.900 ;
      LAYER met1 ;
        RECT 71.050 11.550 79.100 11.900 ;
      LAYER met1 ;
        RECT 79.100 11.550 80.850 13.650 ;
      LAYER met1 ;
        RECT 80.850 11.550 83.300 13.650 ;
      LAYER met1 ;
        RECT 83.300 11.550 85.050 18.200 ;
      LAYER met1 ;
        RECT 85.050 13.650 86.100 18.200 ;
      LAYER met1 ;
        RECT 86.100 15.050 87.850 18.200 ;
      LAYER met1 ;
        RECT 87.850 15.050 93.100 18.200 ;
      LAYER met1 ;
        RECT 93.100 16.450 94.500 19.600 ;
      LAYER met1 ;
        RECT 94.500 19.250 97.650 19.600 ;
      LAYER met1 ;
        RECT 97.650 19.250 98.350 19.600 ;
      LAYER met1 ;
        RECT 98.350 19.250 109.900 19.600 ;
        RECT 94.500 18.900 97.300 19.250 ;
      LAYER met1 ;
        RECT 97.300 18.900 98.700 19.250 ;
      LAYER met1 ;
        RECT 98.700 18.900 109.900 19.250 ;
        RECT 94.500 18.550 96.950 18.900 ;
      LAYER met1 ;
        RECT 96.950 18.550 99.050 18.900 ;
      LAYER met1 ;
        RECT 94.500 18.200 96.600 18.550 ;
      LAYER met1 ;
        RECT 96.600 18.200 99.050 18.550 ;
      LAYER met1 ;
        RECT 99.050 18.200 109.900 18.900 ;
        RECT 94.500 17.850 96.250 18.200 ;
      LAYER met1 ;
        RECT 96.250 17.850 98.700 18.200 ;
      LAYER met1 ;
        RECT 98.700 17.850 109.900 18.200 ;
        RECT 94.500 17.500 95.900 17.850 ;
      LAYER met1 ;
        RECT 95.900 17.500 98.350 17.850 ;
      LAYER met1 ;
        RECT 98.350 17.500 109.900 17.850 ;
        RECT 94.500 17.150 95.550 17.500 ;
      LAYER met1 ;
        RECT 95.550 17.150 98.000 17.500 ;
      LAYER met1 ;
        RECT 98.000 17.150 109.900 17.500 ;
        RECT 94.500 16.450 95.200 17.150 ;
      LAYER met1 ;
        RECT 95.200 16.800 97.650 17.150 ;
      LAYER met1 ;
        RECT 97.650 16.800 109.900 17.150 ;
      LAYER met1 ;
        RECT 95.200 16.450 97.300 16.800 ;
      LAYER met1 ;
        RECT 97.300 16.450 109.900 16.800 ;
      LAYER met1 ;
        RECT 93.100 16.100 96.950 16.450 ;
      LAYER met1 ;
        RECT 96.950 16.100 109.900 16.450 ;
      LAYER met1 ;
        RECT 93.100 15.750 96.600 16.100 ;
      LAYER met1 ;
        RECT 96.600 15.750 109.900 16.100 ;
      LAYER met1 ;
        RECT 93.100 15.400 96.250 15.750 ;
      LAYER met1 ;
        RECT 96.250 15.400 109.900 15.750 ;
      LAYER met1 ;
        RECT 93.100 15.050 95.900 15.400 ;
      LAYER met1 ;
        RECT 95.900 15.050 109.900 15.400 ;
      LAYER met1 ;
        RECT 86.100 13.650 92.050 15.050 ;
      LAYER met1 ;
        RECT 85.050 13.300 90.300 13.650 ;
      LAYER met1 ;
        RECT 90.300 13.300 92.050 13.650 ;
      LAYER met1 ;
        RECT 85.050 11.550 90.650 13.300 ;
      LAYER met1 ;
        RECT 90.650 11.550 92.050 13.300 ;
      LAYER met1 ;
        RECT 64.750 11.200 68.250 11.550 ;
      LAYER met1 ;
        RECT 68.250 11.200 70.350 11.550 ;
      LAYER met1 ;
        RECT 70.350 11.200 79.100 11.550 ;
        RECT 24.500 10.850 29.750 11.200 ;
      LAYER met1 ;
        RECT 29.750 10.850 31.850 11.200 ;
      LAYER met1 ;
        RECT 31.850 10.850 33.600 11.200 ;
      LAYER met1 ;
        RECT 33.600 10.850 35.700 11.200 ;
      LAYER met1 ;
        RECT 35.700 10.850 79.100 11.200 ;
        RECT 19.600 10.500 20.300 10.850 ;
      LAYER met1 ;
        RECT 20.300 10.500 26.600 10.850 ;
      LAYER met1 ;
        RECT 26.600 10.500 30.100 10.850 ;
      LAYER met1 ;
        RECT 30.100 10.500 32.200 10.850 ;
      LAYER met1 ;
        RECT 32.200 10.500 33.250 10.850 ;
      LAYER met1 ;
        RECT 33.250 10.500 35.350 10.850 ;
      LAYER met1 ;
        RECT 35.350 10.500 79.100 10.850 ;
        RECT 19.600 10.150 19.950 10.500 ;
      LAYER met1 ;
        RECT 19.950 10.150 26.600 10.500 ;
      LAYER met1 ;
        RECT 26.600 10.150 30.450 10.500 ;
      LAYER met1 ;
        RECT 30.450 10.150 35.000 10.500 ;
      LAYER met1 ;
        RECT 35.000 10.150 79.100 10.500 ;
        RECT 19.600 9.800 20.300 10.150 ;
      LAYER met1 ;
        RECT 20.300 9.800 26.250 10.150 ;
      LAYER met1 ;
        RECT 26.250 9.800 31.150 10.150 ;
      LAYER met1 ;
        RECT 31.150 9.800 34.300 10.150 ;
      LAYER met1 ;
        RECT 34.300 9.800 79.100 10.150 ;
      LAYER met1 ;
        RECT 79.100 9.800 85.050 11.550 ;
      LAYER met1 ;
        RECT 85.050 9.800 86.100 11.550 ;
      LAYER met1 ;
        RECT 86.100 9.800 92.050 11.550 ;
      LAYER met1 ;
        RECT 92.050 9.800 93.100 15.050 ;
      LAYER met1 ;
        RECT 93.100 14.700 95.550 15.050 ;
      LAYER met1 ;
        RECT 95.550 14.700 109.900 15.050 ;
      LAYER met1 ;
        RECT 93.100 14.350 95.900 14.700 ;
      LAYER met1 ;
        RECT 95.900 14.350 109.900 14.700 ;
      LAYER met1 ;
        RECT 93.100 14.000 96.250 14.350 ;
      LAYER met1 ;
        RECT 96.250 14.000 109.900 14.350 ;
      LAYER met1 ;
        RECT 93.100 13.650 96.600 14.000 ;
      LAYER met1 ;
        RECT 96.600 13.650 109.900 14.000 ;
      LAYER met1 ;
        RECT 93.100 13.300 96.950 13.650 ;
      LAYER met1 ;
        RECT 96.950 13.300 109.900 13.650 ;
      LAYER met1 ;
        RECT 93.100 9.800 94.500 13.300 ;
      LAYER met1 ;
        RECT 94.500 12.950 94.850 13.300 ;
      LAYER met1 ;
        RECT 94.850 12.950 97.300 13.300 ;
      LAYER met1 ;
        RECT 97.300 12.950 109.900 13.300 ;
        RECT 94.500 12.600 95.200 12.950 ;
      LAYER met1 ;
        RECT 95.200 12.600 97.650 12.950 ;
      LAYER met1 ;
        RECT 94.500 12.250 95.550 12.600 ;
      LAYER met1 ;
        RECT 95.550 12.250 97.650 12.600 ;
      LAYER met1 ;
        RECT 97.650 12.250 109.900 12.950 ;
        RECT 94.500 11.900 95.900 12.250 ;
      LAYER met1 ;
        RECT 95.900 11.900 98.000 12.250 ;
      LAYER met1 ;
        RECT 98.000 11.900 109.900 12.250 ;
        RECT 94.500 11.550 96.250 11.900 ;
      LAYER met1 ;
        RECT 96.250 11.550 98.350 11.900 ;
      LAYER met1 ;
        RECT 98.350 11.550 109.900 11.900 ;
        RECT 94.500 11.200 96.600 11.550 ;
      LAYER met1 ;
        RECT 96.600 11.200 98.700 11.550 ;
      LAYER met1 ;
        RECT 98.700 11.200 109.900 11.550 ;
        RECT 94.500 10.850 96.950 11.200 ;
      LAYER met1 ;
        RECT 96.950 10.850 99.050 11.200 ;
      LAYER met1 ;
        RECT 94.500 10.500 97.300 10.850 ;
      LAYER met1 ;
        RECT 97.300 10.500 99.050 10.850 ;
      LAYER met1 ;
        RECT 99.050 10.500 109.900 11.200 ;
        RECT 94.500 10.150 97.650 10.500 ;
      LAYER met1 ;
        RECT 97.650 10.150 98.700 10.500 ;
      LAYER met1 ;
        RECT 98.700 10.150 109.900 10.500 ;
        RECT 94.500 9.800 98.000 10.150 ;
      LAYER met1 ;
        RECT 98.000 9.800 98.350 10.150 ;
      LAYER met1 ;
        RECT 98.350 9.800 109.900 10.150 ;
        RECT 19.600 9.100 109.900 9.800 ;
      LAYER met1 ;
        RECT 0.350 7.350 2.100 7.700 ;
      LAYER met1 ;
        RECT 0.000 6.300 0.700 7.350 ;
      LAYER met1 ;
        RECT 0.700 7.000 2.100 7.350 ;
      LAYER met1 ;
        RECT 2.100 7.000 5.950 7.700 ;
      LAYER met1 ;
        RECT 5.950 7.000 8.750 8.750 ;
      LAYER met1 ;
        RECT 8.750 7.000 10.500 8.750 ;
      LAYER met1 ;
        RECT 0.700 6.300 2.450 7.000 ;
      LAYER met1 ;
        RECT 2.450 6.300 10.500 7.000 ;
        RECT 0.000 5.600 1.050 6.300 ;
      LAYER met1 ;
        RECT 1.050 5.600 2.800 6.300 ;
      LAYER met1 ;
        RECT 2.800 5.600 10.500 6.300 ;
        RECT 0.000 5.250 1.400 5.600 ;
      LAYER met1 ;
        RECT 1.400 5.250 3.150 5.600 ;
      LAYER met1 ;
        RECT 3.150 5.250 10.500 5.600 ;
        RECT 0.000 4.550 1.750 5.250 ;
      LAYER met1 ;
        RECT 1.750 4.900 3.500 5.250 ;
      LAYER met1 ;
        RECT 3.500 4.900 10.500 5.250 ;
      LAYER met1 ;
        RECT 1.750 4.550 3.850 4.900 ;
      LAYER met1 ;
        RECT 3.850 4.550 10.500 4.900 ;
        RECT 0.000 4.200 2.100 4.550 ;
      LAYER met1 ;
        RECT 2.100 4.200 4.200 4.550 ;
      LAYER met1 ;
        RECT 4.200 4.200 10.500 4.550 ;
        RECT 0.000 3.850 2.450 4.200 ;
      LAYER met1 ;
        RECT 2.450 3.850 4.550 4.200 ;
      LAYER met1 ;
        RECT 4.550 3.850 10.500 4.200 ;
        RECT 0.000 3.500 2.800 3.850 ;
      LAYER met1 ;
        RECT 2.800 3.500 4.900 3.850 ;
      LAYER met1 ;
        RECT 4.900 3.500 10.500 3.850 ;
        RECT 0.000 3.150 3.150 3.500 ;
      LAYER met1 ;
        RECT 3.150 3.150 5.600 3.500 ;
      LAYER met1 ;
        RECT 5.600 3.150 10.500 3.500 ;
        RECT 0.000 2.800 3.500 3.150 ;
      LAYER met1 ;
        RECT 3.500 2.800 6.300 3.150 ;
      LAYER met1 ;
        RECT 6.300 2.800 10.500 3.150 ;
        RECT 0.000 2.450 3.850 2.800 ;
      LAYER met1 ;
        RECT 3.850 2.450 7.000 2.800 ;
      LAYER met1 ;
        RECT 7.000 2.450 10.500 2.800 ;
        RECT 0.000 2.100 4.550 2.450 ;
      LAYER met1 ;
        RECT 4.550 2.100 8.400 2.450 ;
      LAYER met1 ;
        RECT 8.400 2.100 10.500 2.450 ;
      LAYER met1 ;
        RECT 10.500 2.100 13.300 8.750 ;
      LAYER met1 ;
        RECT 13.300 8.050 17.850 8.750 ;
      LAYER met1 ;
        RECT 17.850 8.050 19.250 9.100 ;
      LAYER met1 ;
        RECT 19.250 8.050 109.900 9.100 ;
        RECT 13.300 7.000 17.500 8.050 ;
      LAYER met1 ;
        RECT 17.500 7.700 19.250 8.050 ;
      LAYER met1 ;
        RECT 19.250 7.700 40.600 8.050 ;
      LAYER met1 ;
        RECT 17.500 7.000 18.900 7.700 ;
      LAYER met1 ;
        RECT 18.900 7.350 40.600 7.700 ;
        RECT 18.900 7.000 20.300 7.350 ;
      LAYER met1 ;
        RECT 20.300 7.000 22.400 7.350 ;
      LAYER met1 ;
        RECT 22.400 7.000 25.200 7.350 ;
      LAYER met1 ;
        RECT 25.200 7.000 26.600 7.350 ;
      LAYER met1 ;
        RECT 26.600 7.000 29.050 7.350 ;
      LAYER met1 ;
        RECT 29.050 7.000 30.800 7.350 ;
      LAYER met1 ;
        RECT 30.800 7.000 32.900 7.350 ;
        RECT 13.300 6.300 17.150 7.000 ;
      LAYER met1 ;
        RECT 17.150 6.650 18.900 7.000 ;
      LAYER met1 ;
        RECT 18.900 6.650 19.950 7.000 ;
      LAYER met1 ;
        RECT 19.950 6.650 22.750 7.000 ;
      LAYER met1 ;
        RECT 22.750 6.650 24.850 7.000 ;
      LAYER met1 ;
        RECT 24.850 6.650 26.950 7.000 ;
      LAYER met1 ;
        RECT 26.950 6.650 28.350 7.000 ;
      LAYER met1 ;
        RECT 28.350 6.650 31.150 7.000 ;
      LAYER met1 ;
        RECT 31.150 6.650 32.900 7.000 ;
      LAYER met1 ;
        RECT 17.150 6.300 18.550 6.650 ;
      LAYER met1 ;
        RECT 18.550 6.300 19.950 6.650 ;
      LAYER met1 ;
        RECT 19.950 6.300 21.000 6.650 ;
      LAYER met1 ;
        RECT 21.000 6.300 21.700 6.650 ;
      LAYER met1 ;
        RECT 21.700 6.300 23.100 6.650 ;
      LAYER met1 ;
        RECT 13.300 5.950 16.800 6.300 ;
      LAYER met1 ;
        RECT 16.800 5.950 18.550 6.300 ;
      LAYER met1 ;
        RECT 18.550 5.950 22.050 6.300 ;
        RECT 13.300 5.250 16.450 5.950 ;
      LAYER met1 ;
        RECT 16.450 5.250 18.200 5.950 ;
      LAYER met1 ;
        RECT 18.200 5.250 22.050 5.950 ;
      LAYER met1 ;
        RECT 22.050 5.250 23.100 6.300 ;
      LAYER met1 ;
        RECT 23.100 5.950 24.500 6.650 ;
      LAYER met1 ;
        RECT 24.500 6.300 27.300 6.650 ;
      LAYER met1 ;
        RECT 27.300 6.300 28.350 6.650 ;
      LAYER met1 ;
        RECT 28.350 6.300 29.400 6.650 ;
      LAYER met1 ;
        RECT 29.400 6.300 30.100 6.650 ;
      LAYER met1 ;
        RECT 30.100 6.300 31.500 6.650 ;
        RECT 24.500 5.950 25.550 6.300 ;
      LAYER met1 ;
        RECT 25.550 5.950 26.250 6.300 ;
      LAYER met1 ;
        RECT 26.250 5.950 27.300 6.300 ;
      LAYER met1 ;
        RECT 23.100 5.250 24.150 5.950 ;
        RECT 13.300 4.900 16.100 5.250 ;
      LAYER met1 ;
        RECT 16.100 4.900 17.850 5.250 ;
      LAYER met1 ;
        RECT 17.850 4.900 21.700 5.250 ;
        RECT 13.300 4.550 15.750 4.900 ;
      LAYER met1 ;
        RECT 15.750 4.550 17.500 4.900 ;
      LAYER met1 ;
        RECT 17.500 4.550 21.700 4.900 ;
      LAYER met1 ;
        RECT 21.700 4.550 22.750 5.250 ;
      LAYER met1 ;
        RECT 22.750 4.550 24.150 5.250 ;
        RECT 13.300 4.200 15.400 4.550 ;
      LAYER met1 ;
        RECT 15.400 4.200 17.500 4.550 ;
      LAYER met1 ;
        RECT 17.500 4.200 21.350 4.550 ;
      LAYER met1 ;
        RECT 21.350 4.200 22.400 4.550 ;
      LAYER met1 ;
        RECT 22.400 4.200 24.150 4.550 ;
        RECT 13.300 3.850 15.050 4.200 ;
      LAYER met1 ;
        RECT 15.050 3.850 17.150 4.200 ;
      LAYER met1 ;
        RECT 17.150 3.850 21.000 4.200 ;
      LAYER met1 ;
        RECT 21.000 3.850 22.050 4.200 ;
      LAYER met1 ;
        RECT 22.050 3.850 24.150 4.200 ;
        RECT 13.300 3.150 14.350 3.850 ;
      LAYER met1 ;
        RECT 14.350 3.500 16.800 3.850 ;
      LAYER met1 ;
        RECT 16.800 3.500 20.650 3.850 ;
      LAYER met1 ;
        RECT 20.650 3.500 21.700 3.850 ;
      LAYER met1 ;
        RECT 21.700 3.500 24.150 3.850 ;
      LAYER met1 ;
        RECT 24.150 3.500 25.200 5.950 ;
      LAYER met1 ;
        RECT 25.200 4.900 26.600 5.950 ;
      LAYER met1 ;
        RECT 26.600 5.600 27.300 5.950 ;
      LAYER met1 ;
        RECT 27.300 5.600 30.450 6.300 ;
        RECT 25.200 4.200 25.550 4.900 ;
      LAYER met1 ;
        RECT 25.550 4.200 26.250 4.900 ;
      LAYER met1 ;
        RECT 26.250 4.200 26.600 4.900 ;
        RECT 25.200 3.500 26.600 4.200 ;
      LAYER met1 ;
        RECT 26.600 3.500 27.650 5.600 ;
      LAYER met1 ;
        RECT 27.650 4.900 30.450 5.600 ;
      LAYER met1 ;
        RECT 30.450 4.900 31.500 6.300 ;
      LAYER met1 ;
        RECT 31.500 4.900 32.900 6.650 ;
      LAYER met1 ;
        RECT 32.900 6.300 35.700 7.350 ;
      LAYER met1 ;
        RECT 35.700 6.300 40.600 7.350 ;
      LAYER met1 ;
        RECT 40.600 7.000 44.100 8.050 ;
      LAYER met1 ;
        RECT 44.100 7.700 59.500 8.050 ;
      LAYER met1 ;
        RECT 59.500 7.700 59.850 8.050 ;
      LAYER met1 ;
        RECT 59.850 7.700 79.450 8.050 ;
      LAYER met1 ;
        RECT 79.450 7.700 82.950 8.050 ;
      LAYER met1 ;
        RECT 82.950 7.700 109.900 8.050 ;
      LAYER met1 ;
        RECT 40.600 6.650 41.650 7.000 ;
      LAYER met1 ;
        RECT 41.650 6.650 43.050 7.000 ;
      LAYER met1 ;
        RECT 32.900 5.600 33.600 6.300 ;
      LAYER met1 ;
        RECT 33.600 5.600 40.600 6.300 ;
      LAYER met1 ;
        RECT 32.900 5.250 34.650 5.600 ;
      LAYER met1 ;
        RECT 34.650 5.250 40.600 5.600 ;
      LAYER met1 ;
        RECT 40.600 5.250 41.300 6.650 ;
      LAYER met1 ;
        RECT 41.300 5.250 43.050 6.650 ;
      LAYER met1 ;
        RECT 43.050 5.250 44.100 7.000 ;
      LAYER met1 ;
        RECT 44.100 6.650 59.150 7.700 ;
      LAYER met1 ;
        RECT 32.900 4.900 35.350 5.250 ;
      LAYER met1 ;
        RECT 35.350 4.900 40.600 5.250 ;
        RECT 27.650 4.550 30.100 4.900 ;
      LAYER met1 ;
        RECT 30.100 4.550 31.150 4.900 ;
      LAYER met1 ;
        RECT 31.150 4.550 32.900 4.900 ;
      LAYER met1 ;
        RECT 32.900 4.550 35.700 4.900 ;
      LAYER met1 ;
        RECT 27.650 4.200 29.750 4.550 ;
      LAYER met1 ;
        RECT 29.750 4.200 30.800 4.550 ;
      LAYER met1 ;
        RECT 30.800 4.200 34.650 4.550 ;
      LAYER met1 ;
        RECT 34.650 4.200 35.700 4.550 ;
      LAYER met1 ;
        RECT 35.700 4.200 40.600 4.900 ;
      LAYER met1 ;
        RECT 40.600 4.200 44.100 5.250 ;
      LAYER met1 ;
        RECT 27.650 3.850 29.400 4.200 ;
      LAYER met1 ;
        RECT 29.400 3.850 30.450 4.200 ;
      LAYER met1 ;
        RECT 30.450 3.850 35.000 4.200 ;
        RECT 27.650 3.500 29.050 3.850 ;
      LAYER met1 ;
        RECT 29.050 3.500 30.100 3.850 ;
      LAYER met1 ;
        RECT 30.100 3.500 35.000 3.850 ;
      LAYER met1 ;
        RECT 14.350 3.150 16.450 3.500 ;
      LAYER met1 ;
        RECT 16.450 3.150 20.300 3.500 ;
      LAYER met1 ;
        RECT 20.300 3.150 21.350 3.500 ;
      LAYER met1 ;
        RECT 21.350 3.150 24.500 3.500 ;
      LAYER met1 ;
        RECT 24.500 3.150 25.200 3.500 ;
      LAYER met1 ;
        RECT 25.200 3.150 26.250 3.500 ;
        RECT 13.300 2.100 14.000 3.150 ;
      LAYER met1 ;
        RECT 14.000 2.800 16.100 3.150 ;
      LAYER met1 ;
        RECT 16.100 2.800 19.950 3.150 ;
      LAYER met1 ;
        RECT 14.000 2.450 15.750 2.800 ;
      LAYER met1 ;
        RECT 15.750 2.450 19.950 2.800 ;
      LAYER met1 ;
        RECT 14.000 2.100 15.050 2.450 ;
      LAYER met1 ;
        RECT 15.050 2.100 19.950 2.450 ;
      LAYER met1 ;
        RECT 19.950 2.100 23.100 3.150 ;
      LAYER met1 ;
        RECT 23.100 2.450 24.500 3.150 ;
      LAYER met1 ;
        RECT 24.500 2.800 25.550 3.150 ;
      LAYER met1 ;
        RECT 25.550 2.800 26.250 3.150 ;
      LAYER met1 ;
        RECT 26.250 2.800 27.300 3.500 ;
      LAYER met1 ;
        RECT 27.300 3.150 28.700 3.500 ;
      LAYER met1 ;
        RECT 28.700 3.150 29.750 3.500 ;
      LAYER met1 ;
        RECT 29.750 3.150 35.000 3.500 ;
      LAYER met1 ;
        RECT 35.000 3.150 36.050 4.200 ;
      LAYER met1 ;
        RECT 36.050 3.150 40.600 4.200 ;
      LAYER met1 ;
        RECT 40.600 3.850 41.650 4.200 ;
      LAYER met1 ;
        RECT 41.650 3.850 43.050 4.200 ;
        RECT 27.300 2.800 28.350 3.150 ;
      LAYER met1 ;
        RECT 24.500 2.450 26.950 2.800 ;
      LAYER met1 ;
        RECT 23.100 2.100 24.850 2.450 ;
      LAYER met1 ;
        RECT 24.850 2.100 26.950 2.450 ;
      LAYER met1 ;
        RECT 26.950 2.100 28.350 2.800 ;
      LAYER met1 ;
        RECT 28.350 2.100 31.500 3.150 ;
      LAYER met1 ;
        RECT 31.500 2.800 32.900 3.150 ;
      LAYER met1 ;
        RECT 32.900 2.800 33.250 3.150 ;
      LAYER met1 ;
        RECT 33.250 2.800 34.650 3.150 ;
      LAYER met1 ;
        RECT 34.650 2.800 35.700 3.150 ;
      LAYER met1 ;
        RECT 31.500 2.450 32.550 2.800 ;
      LAYER met1 ;
        RECT 32.550 2.450 35.700 2.800 ;
      LAYER met1 ;
        RECT 35.700 2.450 40.600 3.150 ;
      LAYER met1 ;
        RECT 40.600 2.450 41.300 3.850 ;
      LAYER met1 ;
        RECT 41.300 2.450 43.050 3.850 ;
        RECT 31.500 2.100 32.900 2.450 ;
      LAYER met1 ;
        RECT 32.900 2.100 35.350 2.450 ;
      LAYER met1 ;
        RECT 35.350 2.100 40.600 2.450 ;
      LAYER met1 ;
        RECT 40.600 2.100 41.650 2.450 ;
      LAYER met1 ;
        RECT 41.650 2.100 43.050 2.450 ;
      LAYER met1 ;
        RECT 43.050 2.100 44.100 4.200 ;
      LAYER met1 ;
        RECT 44.100 2.100 44.450 6.650 ;
      LAYER met1 ;
        RECT 44.450 6.300 45.500 6.650 ;
      LAYER met1 ;
        RECT 45.500 6.300 47.250 6.650 ;
      LAYER met1 ;
        RECT 44.450 5.600 45.850 6.300 ;
      LAYER met1 ;
        RECT 45.850 5.600 47.250 6.300 ;
      LAYER met1 ;
        RECT 44.450 5.250 46.200 5.600 ;
      LAYER met1 ;
        RECT 46.200 5.250 47.250 5.600 ;
      LAYER met1 ;
        RECT 44.450 4.550 46.550 5.250 ;
      LAYER met1 ;
        RECT 46.550 4.550 47.250 5.250 ;
      LAYER met1 ;
        RECT 44.450 2.100 45.500 4.550 ;
      LAYER met1 ;
        RECT 45.500 3.850 45.850 4.550 ;
      LAYER met1 ;
        RECT 45.850 4.200 46.900 4.550 ;
      LAYER met1 ;
        RECT 46.900 4.200 47.250 4.550 ;
      LAYER met1 ;
        RECT 47.250 4.200 48.300 6.650 ;
        RECT 45.850 3.850 48.300 4.200 ;
      LAYER met1 ;
        RECT 45.500 3.500 46.200 3.850 ;
      LAYER met1 ;
        RECT 46.200 3.500 48.300 3.850 ;
      LAYER met1 ;
        RECT 45.500 2.800 46.550 3.500 ;
      LAYER met1 ;
        RECT 46.550 2.800 48.300 3.500 ;
      LAYER met1 ;
        RECT 45.500 2.450 46.900 2.800 ;
      LAYER met1 ;
        RECT 46.900 2.450 48.300 2.800 ;
      LAYER met1 ;
        RECT 45.500 2.100 47.250 2.450 ;
      LAYER met1 ;
        RECT 47.250 2.100 48.300 2.450 ;
      LAYER met1 ;
        RECT 48.300 2.100 48.650 6.650 ;
      LAYER met1 ;
        RECT 48.650 6.300 49.350 6.650 ;
      LAYER met1 ;
        RECT 49.350 6.300 51.450 6.650 ;
      LAYER met1 ;
        RECT 51.450 6.300 52.150 6.650 ;
        RECT 48.650 5.950 49.700 6.300 ;
      LAYER met1 ;
        RECT 49.700 5.950 51.100 6.300 ;
      LAYER met1 ;
        RECT 48.650 5.250 50.050 5.950 ;
      LAYER met1 ;
        RECT 50.050 5.250 51.100 5.950 ;
      LAYER met1 ;
        RECT 48.650 4.900 50.400 5.250 ;
      LAYER met1 ;
        RECT 50.400 4.900 51.100 5.250 ;
      LAYER met1 ;
        RECT 48.650 4.200 50.750 4.900 ;
      LAYER met1 ;
        RECT 50.750 4.200 51.100 4.900 ;
      LAYER met1 ;
        RECT 51.100 4.200 52.150 6.300 ;
        RECT 48.650 2.100 49.700 4.200 ;
      LAYER met1 ;
        RECT 49.700 3.500 50.050 4.200 ;
      LAYER met1 ;
        RECT 50.050 3.500 52.150 4.200 ;
      LAYER met1 ;
        RECT 49.700 3.150 50.400 3.500 ;
      LAYER met1 ;
        RECT 50.400 3.150 52.150 3.500 ;
      LAYER met1 ;
        RECT 49.700 2.450 50.750 3.150 ;
      LAYER met1 ;
        RECT 50.750 2.450 52.150 3.150 ;
      LAYER met1 ;
        RECT 49.700 2.100 51.100 2.450 ;
      LAYER met1 ;
        RECT 51.100 2.100 52.150 2.450 ;
      LAYER met1 ;
        RECT 52.150 2.100 52.500 6.650 ;
      LAYER met1 ;
        RECT 52.500 6.300 56.000 6.650 ;
      LAYER met1 ;
        RECT 56.000 6.300 59.150 6.650 ;
      LAYER met1 ;
        RECT 52.500 5.600 56.350 6.300 ;
        RECT 52.500 4.550 53.550 5.600 ;
      LAYER met1 ;
        RECT 53.550 4.900 55.300 5.600 ;
      LAYER met1 ;
        RECT 55.300 4.900 56.350 5.600 ;
      LAYER met1 ;
        RECT 53.550 4.550 54.950 4.900 ;
      LAYER met1 ;
        RECT 54.950 4.550 56.350 4.900 ;
        RECT 52.500 3.850 56.350 4.550 ;
      LAYER met1 ;
        RECT 56.350 3.850 59.150 6.300 ;
      LAYER met1 ;
        RECT 52.500 3.500 56.000 3.850 ;
      LAYER met1 ;
        RECT 56.000 3.500 59.150 3.850 ;
      LAYER met1 ;
        RECT 52.500 3.150 53.550 3.500 ;
      LAYER met1 ;
        RECT 53.550 3.150 59.150 3.500 ;
      LAYER met1 ;
        RECT 52.500 2.800 56.000 3.150 ;
      LAYER met1 ;
        RECT 56.000 2.800 59.150 3.150 ;
      LAYER met1 ;
        RECT 52.500 2.100 56.350 2.800 ;
      LAYER met1 ;
        RECT 56.350 2.100 59.150 2.800 ;
      LAYER met1 ;
        RECT 59.150 2.100 60.200 7.700 ;
      LAYER met1 ;
        RECT 60.200 6.650 79.100 7.700 ;
      LAYER met1 ;
        RECT 79.100 7.000 82.950 7.700 ;
      LAYER met1 ;
        RECT 82.950 7.350 107.100 7.700 ;
      LAYER met1 ;
        RECT 107.100 7.350 108.150 7.700 ;
        RECT 79.100 6.650 80.500 7.000 ;
      LAYER met1 ;
        RECT 80.500 6.650 81.900 7.000 ;
        RECT 60.200 3.850 60.550 6.650 ;
      LAYER met1 ;
        RECT 60.550 6.300 64.050 6.650 ;
      LAYER met1 ;
        RECT 64.050 6.300 65.100 6.650 ;
      LAYER met1 ;
        RECT 65.100 6.300 68.250 6.650 ;
        RECT 60.550 5.600 64.400 6.300 ;
      LAYER met1 ;
        RECT 64.400 5.950 64.750 6.300 ;
      LAYER met1 ;
        RECT 64.750 5.950 68.250 6.300 ;
      LAYER met1 ;
        RECT 64.400 5.600 65.100 5.950 ;
      LAYER met1 ;
        RECT 65.100 5.600 68.250 5.950 ;
      LAYER met1 ;
        RECT 68.250 5.600 68.950 6.650 ;
      LAYER met1 ;
        RECT 68.950 5.600 72.100 6.650 ;
        RECT 60.550 4.550 61.600 5.600 ;
      LAYER met1 ;
        RECT 61.600 4.550 67.200 5.600 ;
      LAYER met1 ;
        RECT 67.200 4.550 68.250 5.600 ;
      LAYER met1 ;
        RECT 68.250 4.900 71.400 5.600 ;
      LAYER met1 ;
        RECT 71.400 4.900 72.100 5.600 ;
      LAYER met1 ;
        RECT 68.250 4.550 71.050 4.900 ;
      LAYER met1 ;
        RECT 71.050 4.550 72.100 4.900 ;
        RECT 60.550 3.850 64.400 4.550 ;
      LAYER met1 ;
        RECT 60.200 3.500 63.000 3.850 ;
      LAYER met1 ;
        RECT 63.000 3.500 64.400 3.850 ;
      LAYER met1 ;
        RECT 60.200 3.150 63.350 3.500 ;
      LAYER met1 ;
        RECT 63.350 3.150 64.400 3.500 ;
      LAYER met1 ;
        RECT 60.200 2.800 60.900 3.150 ;
      LAYER met1 ;
        RECT 60.900 2.800 64.400 3.150 ;
      LAYER met1 ;
        RECT 60.200 2.100 60.550 2.800 ;
      LAYER met1 ;
        RECT 60.550 2.100 64.400 2.800 ;
      LAYER met1 ;
        RECT 64.400 2.100 64.750 4.550 ;
      LAYER met1 ;
        RECT 64.750 3.500 68.250 4.550 ;
        RECT 64.750 3.150 65.450 3.500 ;
      LAYER met1 ;
        RECT 65.450 3.150 67.200 3.500 ;
      LAYER met1 ;
        RECT 67.200 3.150 68.250 3.500 ;
        RECT 64.750 2.100 68.250 3.150 ;
      LAYER met1 ;
        RECT 68.250 2.100 68.600 4.550 ;
      LAYER met1 ;
        RECT 68.600 3.500 72.100 4.550 ;
        RECT 68.600 3.150 69.650 3.500 ;
      LAYER met1 ;
        RECT 69.650 3.150 71.400 3.500 ;
      LAYER met1 ;
        RECT 71.400 3.150 72.100 3.500 ;
        RECT 68.600 2.100 72.100 3.150 ;
      LAYER met1 ;
        RECT 72.100 2.100 72.800 6.650 ;
      LAYER met1 ;
        RECT 72.800 5.600 76.300 6.650 ;
      LAYER met1 ;
        RECT 76.300 5.600 79.100 6.650 ;
      LAYER met1 ;
        RECT 72.800 5.250 73.850 5.600 ;
      LAYER met1 ;
        RECT 73.850 5.250 79.100 5.600 ;
      LAYER met1 ;
        RECT 79.100 5.250 80.150 6.650 ;
      LAYER met1 ;
        RECT 80.150 5.250 81.900 6.650 ;
      LAYER met1 ;
        RECT 81.900 5.250 82.950 7.000 ;
      LAYER met1 ;
        RECT 82.950 6.650 107.450 7.350 ;
      LAYER met1 ;
        RECT 107.450 6.650 108.150 7.350 ;
        RECT 72.800 3.150 73.500 5.250 ;
      LAYER met1 ;
        RECT 73.500 3.150 79.100 5.250 ;
      LAYER met1 ;
        RECT 79.100 4.200 82.950 5.250 ;
      LAYER met1 ;
        RECT 82.950 4.200 83.300 6.650 ;
      LAYER met1 ;
        RECT 83.300 5.600 86.800 6.650 ;
        RECT 79.100 3.850 81.900 4.200 ;
      LAYER met1 ;
        RECT 81.900 3.850 83.300 4.200 ;
      LAYER met1 ;
        RECT 72.800 2.100 76.300 3.150 ;
      LAYER met1 ;
        RECT 76.300 2.100 79.100 3.150 ;
      LAYER met1 ;
        RECT 79.100 2.100 80.150 3.850 ;
      LAYER met1 ;
        RECT 80.150 3.500 80.850 3.850 ;
      LAYER met1 ;
        RECT 80.850 3.500 82.250 3.850 ;
      LAYER met1 ;
        RECT 80.150 2.800 81.200 3.500 ;
      LAYER met1 ;
        RECT 81.200 3.150 82.250 3.500 ;
      LAYER met1 ;
        RECT 82.250 3.150 83.300 3.850 ;
      LAYER met1 ;
        RECT 83.300 3.150 84.350 5.600 ;
      LAYER met1 ;
        RECT 84.350 3.150 86.100 5.600 ;
      LAYER met1 ;
        RECT 86.100 3.150 86.800 5.600 ;
      LAYER met1 ;
        RECT 86.800 3.850 87.500 6.650 ;
      LAYER met1 ;
        RECT 87.500 5.600 91.000 6.650 ;
      LAYER met1 ;
        RECT 91.000 5.600 91.700 6.650 ;
      LAYER met1 ;
        RECT 91.700 5.600 94.850 6.650 ;
      LAYER met1 ;
        RECT 94.850 6.300 95.550 6.650 ;
      LAYER met1 ;
        RECT 95.550 6.300 96.250 6.650 ;
        RECT 87.500 4.900 88.200 5.600 ;
      LAYER met1 ;
        RECT 88.200 4.900 93.800 5.600 ;
      LAYER met1 ;
        RECT 87.500 4.550 88.550 4.900 ;
      LAYER met1 ;
        RECT 88.550 4.550 93.800 4.900 ;
      LAYER met1 ;
        RECT 93.800 4.550 94.850 5.600 ;
        RECT 87.500 3.850 91.000 4.550 ;
      LAYER met1 ;
        RECT 86.800 3.150 89.950 3.850 ;
      LAYER met1 ;
        RECT 89.950 3.150 91.000 3.850 ;
        RECT 81.200 2.800 82.600 3.150 ;
      LAYER met1 ;
        RECT 82.600 2.800 83.300 3.150 ;
        RECT 80.150 2.450 81.550 2.800 ;
      LAYER met1 ;
        RECT 81.550 2.450 82.950 2.800 ;
      LAYER met1 ;
        RECT 82.950 2.450 83.300 2.800 ;
        RECT 80.150 2.100 81.900 2.450 ;
      LAYER met1 ;
        RECT 81.900 2.100 82.600 2.450 ;
      LAYER met1 ;
        RECT 82.600 2.100 83.300 2.450 ;
      LAYER met1 ;
        RECT 83.300 2.100 86.800 3.150 ;
      LAYER met1 ;
        RECT 86.800 2.800 87.500 3.150 ;
      LAYER met1 ;
        RECT 87.500 2.800 91.000 3.150 ;
      LAYER met1 ;
        RECT 86.800 2.450 87.150 2.800 ;
      LAYER met1 ;
        RECT 87.150 2.450 91.000 2.800 ;
      LAYER met1 ;
        RECT 86.800 2.100 87.500 2.450 ;
      LAYER met1 ;
        RECT 87.500 2.100 91.000 2.450 ;
      LAYER met1 ;
        RECT 91.000 2.100 91.350 4.550 ;
      LAYER met1 ;
        RECT 91.350 3.500 94.850 4.550 ;
        RECT 91.350 3.150 92.400 3.500 ;
      LAYER met1 ;
        RECT 92.400 3.150 93.800 3.500 ;
      LAYER met1 ;
        RECT 93.800 3.150 94.850 3.500 ;
        RECT 91.350 2.100 94.850 3.150 ;
      LAYER met1 ;
        RECT 94.850 2.100 95.200 6.300 ;
      LAYER met1 ;
        RECT 95.200 3.150 96.250 6.300 ;
      LAYER met1 ;
        RECT 96.250 3.150 99.400 6.650 ;
      LAYER met1 ;
        RECT 95.200 2.800 98.700 3.150 ;
      LAYER met1 ;
        RECT 98.700 2.800 99.400 3.150 ;
      LAYER met1 ;
        RECT 95.200 2.100 99.050 2.800 ;
      LAYER met1 ;
        RECT 99.050 2.100 99.400 2.800 ;
      LAYER met1 ;
        RECT 99.400 2.100 100.100 6.650 ;
      LAYER met1 ;
        RECT 100.100 6.300 100.800 6.650 ;
      LAYER met1 ;
        RECT 100.800 6.300 101.500 6.650 ;
      LAYER met1 ;
        RECT 101.500 6.300 103.250 6.650 ;
        RECT 100.100 2.100 100.450 6.300 ;
      LAYER met1 ;
        RECT 100.450 5.950 101.850 6.300 ;
      LAYER met1 ;
        RECT 101.850 5.950 103.250 6.300 ;
      LAYER met1 ;
        RECT 100.450 5.250 102.200 5.950 ;
      LAYER met1 ;
        RECT 102.200 5.250 103.250 5.950 ;
      LAYER met1 ;
        RECT 100.450 4.900 102.550 5.250 ;
      LAYER met1 ;
        RECT 102.550 4.900 103.250 5.250 ;
      LAYER met1 ;
        RECT 100.450 4.550 102.900 4.900 ;
        RECT 100.450 2.100 101.500 4.550 ;
      LAYER met1 ;
        RECT 101.500 4.200 101.850 4.550 ;
      LAYER met1 ;
        RECT 101.850 4.200 102.900 4.550 ;
      LAYER met1 ;
        RECT 102.900 4.200 103.250 4.900 ;
      LAYER met1 ;
        RECT 103.250 4.200 104.300 6.650 ;
      LAYER met1 ;
        RECT 101.500 3.500 102.200 4.200 ;
      LAYER met1 ;
        RECT 102.200 3.500 104.300 4.200 ;
      LAYER met1 ;
        RECT 101.500 3.150 102.550 3.500 ;
      LAYER met1 ;
        RECT 102.550 3.150 104.300 3.500 ;
      LAYER met1 ;
        RECT 101.500 2.450 102.900 3.150 ;
      LAYER met1 ;
        RECT 102.900 2.450 104.300 3.150 ;
      LAYER met1 ;
        RECT 101.500 2.100 103.250 2.450 ;
      LAYER met1 ;
        RECT 103.250 2.100 104.300 2.450 ;
      LAYER met1 ;
        RECT 104.300 2.100 104.650 6.650 ;
      LAYER met1 ;
        RECT 104.650 5.600 108.150 6.650 ;
        RECT 104.650 3.150 105.700 5.600 ;
      LAYER met1 ;
        RECT 105.700 5.250 107.100 5.600 ;
      LAYER met1 ;
        RECT 107.100 5.250 108.150 5.600 ;
      LAYER met1 ;
        RECT 105.700 3.150 107.450 5.250 ;
      LAYER met1 ;
        RECT 107.450 3.150 108.150 5.250 ;
        RECT 104.650 2.100 108.150 3.150 ;
      LAYER met1 ;
        RECT 108.150 2.100 109.900 7.700 ;
        RECT 0.000 1.750 4.900 2.100 ;
      LAYER met1 ;
        RECT 4.900 1.750 13.300 2.100 ;
      LAYER met1 ;
        RECT 13.300 1.750 14.350 2.100 ;
      LAYER met1 ;
        RECT 14.350 1.750 14.700 2.100 ;
      LAYER met1 ;
        RECT 14.700 1.750 109.900 2.100 ;
        RECT 0.000 1.400 5.600 1.750 ;
      LAYER met1 ;
        RECT 5.600 1.400 13.300 1.750 ;
      LAYER met1 ;
        RECT 13.300 1.400 109.900 1.750 ;
        RECT 0.000 1.050 6.650 1.400 ;
      LAYER met1 ;
        RECT 6.650 1.050 12.950 1.400 ;
      LAYER met1 ;
        RECT 12.950 1.050 109.900 1.400 ;
        RECT 0.000 0.700 7.700 1.050 ;
      LAYER met1 ;
        RECT 7.700 0.700 11.900 1.050 ;
      LAYER met1 ;
        RECT 11.900 0.700 109.900 1.050 ;
        RECT 0.000 0.000 109.900 0.700 ;
  END
END my_logo
END LIBRARY

