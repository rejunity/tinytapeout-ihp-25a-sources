module ROM (
    input clk,
    input [6:0] address,    // 5-bit address input
    output reg [47:0] data  // 4 bit address + 8 bit data
);

always @(posedge clk) begin
    data <=
           // Instructions for setting up LED Driver.
           (address == 7'b0000000) ? {12'b101000001111, 12'b101000001111, 12'b101000001111, 12'b101000001111} :
           (address == 7'b0000001) ? {12'b110000000001, 12'b110000000001, 12'b110000000001, 12'b110000000001} :
           (address == 7'b0000010) ? {12'b101100001111, 12'b101100001111, 12'b101100001111, 12'b101100001111} :
           (address == 7'b0000011) ? {12'b100100000000, 12'b100100000000, 12'b100100000000, 12'b100100000000} :
           // Bitmaps, each address corresponding to 32 LEDs.
           (address == 7'b0000100) ? {12'b000100000000, 12'b000100010111, 12'b000100000000, 12'b000100000000} :
           (address == 7'b0000101) ? {12'b001000000000, 12'b001011010110, 12'b001000000000, 12'b001000000000} :
           (address == 7'b0000110) ? {12'b001100000111, 12'b001111110100, 12'b001111110000, 12'b001100100000} :
           (address == 7'b0000111) ? {12'b010000011111, 12'b010011111000, 12'b010010000000, 12'b010000100000} :
           (address == 7'b0001000) ? {12'b010101111111, 12'b010111110000, 12'b010111000111, 12'b010110111100} :
           (address == 7'b0001001) ? {12'b011001111111, 12'b011011110000, 12'b011010000000, 12'b011000100000} :
           (address == 7'b0001010) ? {12'b011101111000, 12'b011111010000, 12'b011111110000, 12'b011100100000} :
           (address == 7'b0001011) ? {12'b100000110000, 12'b100000010000, 12'b100000000000, 12'b100000000000} :
           // Bitmaps, each address corresponding to 32 LEDs.
           (address == 7'b0001100) ? {12'b000100000000, 12'b000100000000, 12'b000100000000, 12'b000100000000} :
           (address == 7'b0001101) ? {12'b001000111110, 12'b001001111111, 12'b001001101111, 12'b001000000000} :
           (address == 7'b0001110) ? {12'b001100111110, 12'b001100000011, 12'b001101101111, 12'b001101000001} :
           (address == 7'b0001111) ? {12'b010001001001, 12'b010001111111, 12'b010001101011, 12'b010001111111} :
           (address == 7'b0010000) ? {12'b010101001001, 12'b010101111111, 12'b010101101011, 12'b010101111111} :
           (address == 7'b0010001) ? {12'b011001111111, 12'b011000000011, 12'b011001111011, 12'b011001000001} :
           (address == 7'b0010010) ? {12'b011101111111, 12'b011101111111, 12'b011101111011, 12'b011100000000} :
                                     {12'b100000000000, 12'b100000000000, 12'b100000000000, 12'b100000000000};
end

endmodule
