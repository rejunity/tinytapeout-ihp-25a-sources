module id_rom (
  input wire [7:0] addr,
  output wire [3:0] data
);

  reg [3:0] mem[255:0];
  initial begin
    mem[0] = 4'h0;
    mem[1] = 4'h0;
    mem[2] = 4'h0;
    mem[3] = 4'h0;
    mem[4] = 4'h0;
    mem[5] = 4'h0;
    mem[6] = 4'h0;
    mem[7] = 4'h0;
    mem[8] = 4'h0;
    mem[9] = 4'h0;
    mem[10] = 4'h0;
    mem[11] = 4'h0;
    mem[12] = 4'h0;
    mem[13] = 4'h0;
    mem[14] = 4'h0;
    mem[15] = 4'h0;
    mem[16] = 4'h0;
    mem[17] = 4'h3;
    mem[18] = 4'hC;
    mem[19] = 4'h0;
    mem[20] = 4'h0;
    mem[21] = 4'h0;
    mem[22] = 4'h0;
    mem[23] = 4'h0;
    mem[24] = 4'h0;
    mem[25] = 4'h0;
    mem[26] = 4'h0;
    mem[27] = 4'h0;
    mem[28] = 4'h0;
    mem[29] = 4'h0;
    mem[30] = 4'h0;
    mem[31] = 4'h0;
    mem[32] = 4'h0;
    mem[33] = 4'h4;
    mem[34] = 4'h2;
    mem[35] = 4'h0;
    mem[36] = 4'h0;
    mem[37] = 4'h0;
    mem[38] = 4'h0;
    mem[39] = 4'h0;
    mem[40] = 4'h0;
    mem[41] = 4'h0;
    mem[42] = 4'h0;
    mem[43] = 4'h0;
    mem[44] = 4'h0;
    mem[45] = 4'h0;
    mem[46] = 4'h0;
    mem[47] = 4'h0;
    mem[48] = 4'h0;
    mem[49] = 4'h4;
    mem[50] = 4'h2;
    mem[51] = 4'h0;
    mem[52] = 4'h0;
    mem[53] = 4'h0;
    mem[54] = 4'h0;
    mem[55] = 4'h0;
    mem[56] = 4'h0;
    mem[57] = 4'h0;
    mem[58] = 4'h0;
    mem[59] = 4'h0;
    mem[60] = 4'h0;
    mem[61] = 4'h0;
    mem[62] = 4'h0;
    mem[63] = 4'h0;
    mem[64] = 4'h0;
    mem[65] = 4'h8;
    mem[66] = 4'h1;
    mem[67] = 4'h1;
    mem[68] = 4'hD;
    mem[69] = 4'hD;
    mem[70] = 4'h9;
    mem[71] = 4'h4;
    mem[72] = 4'h7;
    mem[73] = 4'h2;
    mem[74] = 4'h6;
    mem[75] = 4'h7;
    mem[76] = 4'h2;
    mem[77] = 4'h5;
    mem[78] = 4'h7;
    mem[79] = 4'h0;
    mem[80] = 4'h0;
    mem[81] = 4'hF;
    mem[82] = 4'h1;
    mem[83] = 4'h0;
    mem[84] = 4'h8;
    mem[85] = 4'h9;
    mem[86] = 4'h5;
    mem[87] = 4'h4;
    mem[88] = 4'h2;
    mem[89] = 4'h5;
    mem[90] = 4'h5;
    mem[91] = 4'h4;
    mem[92] = 4'h5;
    mem[93] = 4'h5;
    mem[94] = 4'h2;
    mem[95] = 4'h0;
    mem[96] = 4'h0;
    mem[97] = 4'h2;
    mem[98] = 4'h1;
    mem[99] = 4'h0;
    mem[100] = 4'h8;
    mem[101] = 4'h9;
    mem[102] = 4'h5;
    mem[103] = 4'h4;
    mem[104] = 4'h2;
    mem[105] = 4'h5;
    mem[106] = 4'h5;
    mem[107] = 4'h4;
    mem[108] = 4'h5;
    mem[109] = 4'h5;
    mem[110] = 4'h2;
    mem[111] = 4'h0;
    mem[112] = 4'h0;
    mem[113] = 4'hA;
    mem[114] = 4'h1;
    mem[115] = 4'h0;
    mem[116] = 4'h8;
    mem[117] = 4'h9;
    mem[118] = 4'h4;
    mem[119] = 4'h8;
    mem[120] = 4'h2;
    mem[121] = 4'h5;
    mem[122] = 4'h5;
    mem[123] = 4'h6;
    mem[124] = 4'h5;
    mem[125] = 4'h5;
    mem[126] = 4'h2;
    mem[127] = 4'h0;
    mem[128] = 4'h0;
    mem[129] = 4'hB;
    mem[130] = 4'hD;
    mem[131] = 4'h0;
    mem[132] = 4'h8;
    mem[133] = 4'h9;
    mem[134] = 4'h4;
    mem[135] = 4'h8;
    mem[136] = 4'h2;
    mem[137] = 4'h7;
    mem[138] = 4'h6;
    mem[139] = 4'h4;
    mem[140] = 4'h5;
    mem[141] = 4'h5;
    mem[142] = 4'h2;
    mem[143] = 4'h0;
    mem[144] = 4'h0;
    mem[145] = 4'hA;
    mem[146] = 4'h9;
    mem[147] = 4'h0;
    mem[148] = 4'h8;
    mem[149] = 4'h9;
    mem[150] = 4'h4;
    mem[151] = 4'h8;
    mem[152] = 4'h2;
    mem[153] = 4'h5;
    mem[154] = 4'h4;
    mem[155] = 4'h4;
    mem[156] = 4'h5;
    mem[157] = 4'h5;
    mem[158] = 4'h2;
    mem[159] = 4'h0;
    mem[160] = 4'h0;
    mem[161] = 4'hA;
    mem[162] = 4'h9;
    mem[163] = 4'h0;
    mem[164] = 4'h8;
    mem[165] = 4'h9;
    mem[166] = 4'h4;
    mem[167] = 4'h8;
    mem[168] = 4'h2;
    mem[169] = 4'h5;
    mem[170] = 4'h4;
    mem[171] = 4'h4;
    mem[172] = 4'h5;
    mem[173] = 4'h5;
    mem[174] = 4'h2;
    mem[175] = 4'h0;
    mem[176] = 4'h0;
    mem[177] = 4'h8;
    mem[178] = 4'h9;
    mem[179] = 4'h0;
    mem[180] = 4'h9;
    mem[181] = 4'hD;
    mem[182] = 4'h4;
    mem[183] = 4'h8;
    mem[184] = 4'h2;
    mem[185] = 4'h5;
    mem[186] = 4'h4;
    mem[187] = 4'h7;
    mem[188] = 4'h2;
    mem[189] = 4'h2;
    mem[190] = 4'h2;
    mem[191] = 4'h0;
    mem[192] = 4'h0;
    mem[193] = 4'h4;
    mem[194] = 4'hA;
    mem[195] = 4'h0;
    mem[196] = 4'h0;
    mem[197] = 4'h0;
    mem[198] = 4'h0;
    mem[199] = 4'h0;
    mem[200] = 4'h0;
    mem[201] = 4'h0;
    mem[202] = 4'h0;
    mem[203] = 4'h0;
    mem[204] = 4'h0;
    mem[205] = 4'h0;
    mem[206] = 4'h0;
    mem[207] = 4'h0;
    mem[208] = 4'h0;
    mem[209] = 4'h4;
    mem[210] = 4'hA;
    mem[211] = 4'h0;
    mem[212] = 4'h0;
    mem[213] = 4'h0;
    mem[214] = 4'h0;
    mem[215] = 4'h0;
    mem[216] = 4'h0;
    mem[217] = 4'h0;
    mem[218] = 4'h0;
    mem[219] = 4'h0;
    mem[220] = 4'h0;
    mem[221] = 4'h0;
    mem[222] = 4'h0;
    mem[223] = 4'h0;
    mem[224] = 4'h0;
    mem[225] = 4'h3;
    mem[226] = 4'h8;
    mem[227] = 4'h0;
    mem[228] = 4'h0;
    mem[229] = 4'h0;
    mem[230] = 4'h0;
    mem[231] = 4'h0;
    mem[232] = 4'h0;
    mem[233] = 4'h0;
    mem[234] = 4'h0;
    mem[235] = 4'h0;
    mem[236] = 4'h0;
    mem[237] = 4'h0;
    mem[238] = 4'h0;
    mem[239] = 4'h0;
    mem[240] = 4'h0;
    mem[241] = 4'h0;
    mem[242] = 4'h0;
    mem[243] = 4'h0;
    mem[244] = 4'h0;
    mem[245] = 4'h0;
    mem[246] = 4'h0;
    mem[247] = 4'h0;
    mem[248] = 4'h0;
    mem[249] = 4'h0;
    mem[250] = 4'h0;
    mem[251] = 4'h0;
    mem[252] = 4'h0;
    mem[253] = 4'h0;
    mem[254] = 4'h0;
    mem[255] = 4'h0;
  end

  assign data = mem[addr];

endmodule
